-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
	--bootloader sdram
000000 => x"EA000006",
000001 => x"EAFFFFFE",
000002 => x"EAFFFFFE",
000003 => x"EAFFFFFE",
000004 => x"EAFFFFFE",
000005 => x"E1A00000",
000006 => x"EAFFFFFE",
000007 => x"EAFFFFFE",
000008 => x"E59F0040",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA018",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"E1A04000",
000023 => x"E3A00000",
000024 => x"E1A0F004",
000025 => x"EAFFFFFE",
000026 => x"00002000",
000027 => x"00010780",
000028 => x"E3E03A0F",
000029 => x"E5131FFB",
000030 => x"E20020FF",
000031 => x"E3A00001",
000032 => x"E0010210",
000033 => x"E1A0F00E",
000034 => x"E3E03A0F",
000035 => x"E5130FFB",
000036 => x"E1A0F00E",
000037 => x"E3E01A0F",
000038 => x"E5113FFF",
000039 => x"E20000FF",
000040 => x"E3A02001",
000041 => x"E1833012",
000042 => x"E5013FFF",
000043 => x"E1A0F00E",
000044 => x"E20000FF",
000045 => x"E3A02001",
000046 => x"E1A02012",
000047 => x"E3E01A0F",
000048 => x"E5113FFF",
000049 => x"E1E02002",
000050 => x"E0033002",
000051 => x"E5013FFF",
000052 => x"E1A0F00E",
000053 => x"E3E01A0F",
000054 => x"E5113FFF",
000055 => x"E20000FF",
000056 => x"E3A02001",
000057 => x"E0233012",
000058 => x"E5013FFF",
000059 => x"E1A0F00E",
000060 => x"E3E03A0F",
000061 => x"E5030FFF",
000062 => x"E1A0F00E",
000063 => x"E3E02A0F",
000064 => x"E5123EFB",
000065 => x"E3130002",
000066 => x"E3E00000",
000067 => x"15120EFF",
000068 => x"E1A0F00E",
000069 => x"E3E02A0F",
000070 => x"E5123EFB",
000071 => x"E3130001",
000072 => x"0AFFFFFC",
000073 => x"E20030FF",
000074 => x"E5023EFF",
000075 => x"E1A0F00E",
000076 => x"E20000FF",
000077 => x"E3500001",
000078 => x"E3812B01",
000079 => x"03E03A0F",
000080 => x"E3811B09",
000081 => x"13E03A0F",
000082 => x"05031FCF",
000083 => x"15032FCF",
000084 => x"E1A0F00E",
000085 => x"E3E03A0F",
000086 => x"E5030FCB",
000087 => x"E1A0F00E",
000088 => x"E3E02A0F",
000089 => x"E5123FCF",
000090 => x"E3130C01",
000091 => x"1AFFFFFC",
000092 => x"E5020FBF",
000093 => x"E5123FCF",
000094 => x"E3833C01",
000095 => x"E5023FCF",
000096 => x"E3E02A0F",
000097 => x"E5123FCF",
000098 => x"E3130C01",
000099 => x"1AFFFFFC",
000100 => x"E5120FBF",
000101 => x"E1A0F00E",
000102 => x"E3E01A0F",
000103 => x"E5113FC7",
000104 => x"E20000FF",
000105 => x"E3A02001",
000106 => x"E1833012",
000107 => x"E5013FC7",
000108 => x"E1A0F00E",
000109 => x"E20000FF",
000110 => x"E3A02001",
000111 => x"E1A02012",
000112 => x"E3E01A0F",
000113 => x"E5113FC7",
000114 => x"E1E02002",
000115 => x"E0033002",
000116 => x"E5013FC7",
000117 => x"E1A0F00E",
000118 => x"E3E02A0F",
000119 => x"E5123F97",
000120 => x"E1A01420",
000121 => x"E3C33080",
000122 => x"E5023F97",
000123 => x"E5020F9F",
000124 => x"E5021F9B",
000125 => x"E5123F97",
000126 => x"E3833080",
000127 => x"E5023F97",
000128 => x"E1A0F00E",
000129 => x"E92D4030",
000130 => x"E3A0C090",
000131 => x"E20140FE",
000132 => x"E3E0EA0F",
000133 => x"E5DD500F",
000134 => x"E20000FF",
000135 => x"E50E4F93",
000136 => x"E20110FF",
000137 => x"E50ECFAF",
000138 => x"E1A04002",
000139 => x"E203C0FF",
000140 => x"E51E3FAF",
000141 => x"E3130002",
000142 => x"1AFFFFFC",
000143 => x"E51E3FAF",
000144 => x"E3130080",
000145 => x"13E00000",
000146 => x"18BD8030",
000147 => x"E35C0000",
000148 => x"0A000012",
000149 => x"E24C3001",
000150 => x"E203C0FF",
000151 => x"E35C0001",
000152 => x"01A02424",
000153 => x"03E03A0F",
000154 => x"13E03A0F",
000155 => x"05032F93",
000156 => x"15034F93",
000157 => x"E3E02A0F",
000158 => x"E3A03010",
000159 => x"E5023FAF",
000160 => x"E5123FAF",
000161 => x"E3130002",
000162 => x"1AFFFFFC",
000163 => x"E5123FAF",
000164 => x"E3130080",
000165 => x"0AFFFFEC",
000166 => x"E3E00001",
000167 => x"E8BD8030",
000168 => x"E3500077",
000169 => x"1A00000C",
000170 => x"E3E03A0F",
000171 => x"E3A02050",
000172 => x"E5035F93",
000173 => x"E5032FAF",
000174 => x"E1A02003",
000175 => x"E5123FAF",
000176 => x"E3130002",
000177 => x"1AFFFFFC",
000178 => x"E5123FAF",
000179 => x"E2130080",
000180 => x"08BD8030",
000181 => x"E3E00002",
000182 => x"E8BD8030",
000183 => x"E3500072",
000184 => x"13E00003",
000185 => x"18BD8030",
000186 => x"E3813001",
000187 => x"E3E02A0F",
000188 => x"E3A01090",
000189 => x"E5023F93",
000190 => x"E5021FAF",
000191 => x"E5123FAF",
000192 => x"E3130002",
000193 => x"1AFFFFFC",
000194 => x"E5123FAF",
000195 => x"E3130080",
000196 => x"1AFFFFEF",
000197 => x"E3A03068",
000198 => x"E5023FAF",
000199 => x"E3E00A0F",
000200 => x"E5103FAF",
000201 => x"E3130002",
000202 => x"1AFFFFFC",
000203 => x"E5100F93",
000204 => x"E8BD8030",
000205 => x"E20000FF",
000206 => x"E350000F",
000207 => x"979FF100",
000208 => x"EA00000F",
000209 => x"00010404",
000210 => x"000103FC",
000211 => x"000103F4",
000212 => x"000103EC",
000213 => x"000103E4",
000214 => x"000103DC",
000215 => x"000103D4",
000216 => x"000103CC",
000217 => x"000103C4",
000218 => x"000103BC",
000219 => x"000103B4",
000220 => x"000103AC",
000221 => x"000103A4",
000222 => x"0001039C",
000223 => x"00010394",
000224 => x"0001038C",
000225 => x"E3A00000",
000226 => x"E1A0F00E",
000227 => x"EE1F0F1F",
000228 => x"E1A0F00E",
000229 => x"EE1E0F1E",
000230 => x"E1A0F00E",
000231 => x"EE1D0F1D",
000232 => x"E1A0F00E",
000233 => x"EE1C0F1C",
000234 => x"E1A0F00E",
000235 => x"EE1B0F1B",
000236 => x"E1A0F00E",
000237 => x"EE1A0F1A",
000238 => x"E1A0F00E",
000239 => x"EE190F19",
000240 => x"E1A0F00E",
000241 => x"EE180F18",
000242 => x"E1A0F00E",
000243 => x"EE170F17",
000244 => x"E1A0F00E",
000245 => x"EE160F16",
000246 => x"E1A0F00E",
000247 => x"EE150F15",
000248 => x"E1A0F00E",
000249 => x"EE140F14",
000250 => x"E1A0F00E",
000251 => x"EE130F13",
000252 => x"E1A0F00E",
000253 => x"EE120F12",
000254 => x"E1A0F00E",
000255 => x"EE110F11",
000256 => x"E1A0F00E",
000257 => x"EE100F10",
000258 => x"E1A0F00E",
000259 => x"E20110FF",
000260 => x"E2411006",
000261 => x"E3510007",
000262 => x"979FF101",
000263 => x"EA000008",
000264 => x"00010448",
000265 => x"00010444",
000266 => x"00010444",
000267 => x"00010444",
000268 => x"00010444",
000269 => x"00010450",
000270 => x"00010458",
000271 => x"00010440",
000272 => x"EE0D0F1D",
000273 => x"E1A0F00E",
000274 => x"EE060F16",
000275 => x"E1A0F00E",
000276 => x"EE0B0F1B",
000277 => x"E1A0F00E",
000278 => x"EE0C0F1C",
000279 => x"E1A0F00E",
000280 => x"E92D4010",
000281 => x"E1A04000",
000282 => x"E5D00000",
000283 => x"E3500000",
000284 => x"1A000003",
000285 => x"EA000005",
000286 => x"E5F40001",
000287 => x"E3500000",
000288 => x"0A000002",
000289 => x"EBFFFF22",
000290 => x"E3500000",
000291 => x"CAFFFFF9",
000292 => x"E1A00004",
000293 => x"E8BD8010",
000294 => x"E92D4070",
000295 => x"E2514000",
000296 => x"E1A05000",
000297 => x"E20260FF",
000298 => x"DA00000B",
000299 => x"EBFFFF12",
000300 => x"E3700001",
000301 => x"E20030FF",
000302 => x"0A000005",
000303 => x"E3560001",
000304 => x"E5C53000",
000305 => x"E1A00003",
000306 => x"E2855001",
000307 => x"0A000005",
000308 => x"E2444001",
000309 => x"E3540000",
000310 => x"CAFFFFF3",
000311 => x"E59F300C",
000312 => x"E5C53000",
000313 => x"E8BD8070",
000314 => x"EBFFFF09",
000315 => x"EAFFFFF7",
000316 => x"00011060",
000317 => x"E92D4030",
000318 => x"E2514000",
000319 => x"E1A05000",
000320 => x"D8BD8030",
000321 => x"E4D50001",
000322 => x"EBFFFF01",
000323 => x"E2544001",
000324 => x"1AFFFFFB",
000325 => x"E8BD8030",
000326 => x"E92D4010",
000327 => x"E20240FF",
000328 => x"E3540008",
000329 => x"83A04008",
000330 => x"8A000001",
000331 => x"E3540000",
000332 => x"03A04001",
000333 => x"E1A02001",
000334 => x"E1A0E004",
000335 => x"E1A0310E",
000336 => x"E35E0001",
000337 => x"E2433004",
000338 => x"E1A0C000",
000339 => x"81A0C330",
000340 => x"E24E3001",
000341 => x"E20CC00F",
000342 => x"E203E0FF",
000343 => x"E35C0009",
000344 => x"E28C3030",
000345 => x"828C3037",
000346 => x"E35E0000",
000347 => x"E4C23001",
000348 => x"1AFFFFF1",
000349 => x"E2443001",
000350 => x"E20330FF",
000351 => x"E0813003",
000352 => x"E5C3E001",
000353 => x"E8BD8010",
000354 => x"E92D4010",
000355 => x"E1A04000",
000356 => x"E3540007",
000357 => x"E3A01010",
000358 => x"E3A00001",
000359 => x"9A000001",
000360 => x"E3A00000",
000361 => x"E8BD8010",
000362 => x"EBFFFEE0",
000363 => x"E3A00006",
000364 => x"EBFFFEF8",
000365 => x"E3A00000",
000366 => x"EBFFFEE8",
000367 => x"E1A00584",
000368 => x"E8BD4010",
000369 => x"EAFFFEE5",
000370 => x"E0603280",
000371 => x"E0800103",
000372 => x"E0800100",
000373 => x"E1A00200",
000374 => x"E3500000",
000375 => x"D1A0F00E",
000376 => x"E1A00000",
000377 => x"E2500001",
000378 => x"1AFFFFFC",
000379 => x"E1A0F00E",
000380 => x"E212C0FF",
000381 => x"0A00000B",
000382 => x"E5D02000",
000383 => x"E5D13000",
000384 => x"E1520003",
000385 => x"0A000004",
000386 => x"EA000008",
000387 => x"E5F02001",
000388 => x"E5F13001",
000389 => x"E1520003",
000390 => x"1A000004",
000391 => x"E24C3001",
000392 => x"E213C0FF",
000393 => x"1AFFFFF8",
000394 => x"E3A00001",
000395 => x"E1A0F00E",
000396 => x"E3A00000",
000397 => x"E1A0F00E",
000398 => x"E92D4030",
000399 => x"E1A04081",
000400 => x"E3540000",
000401 => x"E1A05000",
000402 => x"D3A00000",
000403 => x"D8BD8030",
000404 => x"E3A00000",
000405 => x"E1A01000",
000406 => x"E7D12005",
000407 => x"E2423030",
000408 => x"E082C200",
000409 => x"E3530009",
000410 => x"E242E041",
000411 => x"924C0030",
000412 => x"9A000007",
000413 => x"E0823200",
000414 => x"E35E0005",
000415 => x"E242C061",
000416 => x"92430037",
000417 => x"9A000002",
000418 => x"E0823200",
000419 => x"E35C0005",
000420 => x"92430057",
000421 => x"E2811001",
000422 => x"E1510004",
000423 => x"1AFFFFED",
000424 => x"E8BD8030",
000425 => x"E52DE004",
000426 => x"E59F0074",
000427 => x"EBFFFF6B",
000428 => x"E59F0070",
000429 => x"EBFFFF69",
000430 => x"E59F006C",
000431 => x"EBFFFF67",
000432 => x"E59F0068",
000433 => x"EBFFFF65",
000434 => x"E59F0064",
000435 => x"EBFFFF63",
000436 => x"E59F0060",
000437 => x"EBFFFF61",
000438 => x"E59F005C",
000439 => x"EBFFFF5F",
000440 => x"E59F0058",
000441 => x"EBFFFF5D",
000442 => x"E59F0054",
000443 => x"EBFFFF5B",
000444 => x"E59F0050",
000445 => x"EBFFFF59",
000446 => x"E59F004C",
000447 => x"EBFFFF57",
000448 => x"E59F0048",
000449 => x"EBFFFF55",
000450 => x"E59F0044",
000451 => x"EBFFFF53",
000452 => x"E59F0040",
000453 => x"EBFFFF51",
000454 => x"E59F003C",
000455 => x"E49DE004",
000456 => x"EAFFFF4E",
000457 => x"00011064",
000458 => x"000110B0",
000459 => x"000110F8",
000460 => x"00011140",
000461 => x"00011188",
000462 => x"000111D0",
000463 => x"00011218",
000464 => x"00011258",
000465 => x"00011290",
000466 => x"000112B4",
000467 => x"000112FC",
000468 => x"00011368",
000469 => x"000113A0",
000470 => x"00011404",
000471 => x"00011468",
000472 => x"E5D03003",
000473 => x"E5D02002",
000474 => x"E5D01000",
000475 => x"E1833402",
000476 => x"E5D00001",
000477 => x"E1833C01",
000478 => x"E1830800",
000479 => x"E1A0F00E",
000480 => x"E92D47F0",
000481 => x"E3A00000",
000482 => x"E24DD018",
000483 => x"EBFFFE57",
000484 => x"E3A0100D",
000485 => x"E3A000C3",
000486 => x"EBFFFF1B",
000487 => x"E3A00063",
000488 => x"EBFFFE8C",
000489 => x"E3A00006",
000490 => x"EBFFFEE1",
000491 => x"E3A01006",
000492 => x"E3800008",
000493 => x"EBFFFF14",
000494 => x"E3A0000D",
000495 => x"EBFFFEDC",
000496 => x"E1A008A0",
000497 => x"E1E00000",
000498 => x"E200000F",
000499 => x"E3500001",
000500 => x"03A04030",
000501 => x"028D9006",
000502 => x"028DA00F",
000503 => x"0A00001A",
000504 => x"E3500002",
000505 => x"0A000077",
000506 => x"EBFFFFAD",
000507 => x"E28D9006",
000508 => x"E59F07B4",
000509 => x"EBFFFF19",
000510 => x"E1A01009",
000511 => x"E3A02008",
000512 => x"E28D0014",
000513 => x"EBFFFF43",
000514 => x"E1A00009",
000515 => x"EBFFFF13",
000516 => x"E59F0798",
000517 => x"EBFFFF11",
000518 => x"E59F0794",
000519 => x"EBFFFF0F",
000520 => x"E1A01009",
000521 => x"E3A02008",
000522 => x"E3A00301",
000523 => x"EBFFFF39",
000524 => x"E1A00009",
000525 => x"EBFFFF09",
000526 => x"E59F0770",
000527 => x"EBFFFF07",
000528 => x"E28DA00F",
000529 => x"EBFFFE2C",
000530 => x"E1A04000",
000531 => x"E3A0000D",
000532 => x"EBFFFEB7",
000533 => x"E3100801",
000534 => x"03A06001",
000535 => x"03A040A0",
000536 => x"1A00003C",
000537 => x"E3A05000",
000538 => x"E59F0748",
000539 => x"EBFFFEFB",
000540 => x"E1A01004",
000541 => x"E1A02005",
000542 => x"E3A03002",
000543 => x"E3A00072",
000544 => x"E58D5000",
000545 => x"EBFFFE5E",
000546 => x"E1A01004",
000547 => x"E5CD000F",
000548 => x"E3A02001",
000549 => x"E3A03002",
000550 => x"E3A00072",
000551 => x"E58D5000",
000552 => x"EBFFFE57",
000553 => x"E3A02002",
000554 => x"E1A03002",
000555 => x"E5CD0010",
000556 => x"E1A01004",
000557 => x"E3A00072",
000558 => x"E58D5000",
000559 => x"EBFFFE50",
000560 => x"E3A03002",
000561 => x"E5CD0011",
000562 => x"E1A01004",
000563 => x"E3A00072",
000564 => x"E3A02003",
000565 => x"E58D5000",
000566 => x"EBFFFE49",
000567 => x"E5DD300F",
000568 => x"E20000FF",
000569 => x"E3530053",
000570 => x"E5CD0012",
000571 => x"1A000002",
000572 => x"E5DD3010",
000573 => x"E353004D",
000574 => x"0A00006A",
000575 => x"E59F06B8",
000576 => x"EBFFFED6",
000577 => x"E3560000",
000578 => x"0AFFFFCD",
000579 => x"E59F06AC",
000580 => x"EBFFFED2",
000581 => x"E3A0100D",
000582 => x"E3A00000",
000583 => x"EBFFFEBA",
000584 => x"E59F069C",
000585 => x"EBFFFECD",
000586 => x"E3A00006",
000587 => x"EBFFFE80",
000588 => x"E3A01006",
000589 => x"E3C00008",
000590 => x"EBFFFEB3",
000591 => x"E59F0684",
000592 => x"EBFFFEC6",
000593 => x"E3A00301",
000594 => x"EBFFFDC2",
000595 => x"E59F0678",
000596 => x"EBFFFEC2",
000597 => x"EAFFFFFE",
000598 => x"E3540034",
000599 => x"0A000029",
000600 => x"CA00001C",
000601 => x"E3540031",
000602 => x"0A000036",
000603 => x"DA00009B",
000604 => x"E3540032",
000605 => x"0A0000A5",
000606 => x"E3540033",
000607 => x"1A00009B",
000608 => x"E1A00004",
000609 => x"EBFFFDE2",
000610 => x"E59F0640",
000611 => x"EBFFFEB3",
000612 => x"E1A0000A",
000613 => x"E3A01002",
000614 => x"E3A02001",
000615 => x"EBFFFEBD",
000616 => x"E3A01002",
000617 => x"E1A0000A",
000618 => x"EBFFFF22",
000619 => x"E21010FF",
000620 => x"11A04001",
000621 => x"13A06000",
000622 => x"1AFFFFA9",
000623 => x"E59F0610",
000624 => x"EBFFFEA6",
000625 => x"EAFFFF9E",
000626 => x"E3A04033",
000627 => x"E28D9006",
000628 => x"E28DA00F",
000629 => x"EAFFFF9C",
000630 => x"E3540066",
000631 => x"0A00002A",
000632 => x"DA0000B0",
000633 => x"E3540068",
000634 => x"0A000112",
000635 => x"E3540072",
000636 => x"1A00007E",
000637 => x"E1A00004",
000638 => x"EBFFFDC5",
000639 => x"E3A006FF",
000640 => x"E280F20F",
000641 => x"EAFFFFFE",
000642 => x"E1A00004",
000643 => x"EBFFFDC0",
000644 => x"E59F05B8",
000645 => x"EBFFFE91",
000646 => x"E1A0000A",
000647 => x"E3A01002",
000648 => x"E3A02001",
000649 => x"EBFFFE9B",
000650 => x"E1A0000A",
000651 => x"E3A01002",
000652 => x"EBFFFF00",
000653 => x"E21080FF",
000654 => x"1A0000A7",
000655 => x"E59F0594",
000656 => x"EBFFFE86",
000657 => x"EAFFFF7E",
000658 => x"E1A00004",
000659 => x"EBFFFDB0",
000660 => x"E59F0584",
000661 => x"EBFFFE81",
000662 => x"E1A0000A",
000663 => x"E3A01004",
000664 => x"E3A02000",
000665 => x"EBFFFE8B",
000666 => x"E5DD300F",
000667 => x"E3530053",
000668 => x"1A000002",
000669 => x"E5DD3010",
000670 => x"E353004D",
000671 => x"0A0000F1",
000672 => x"E59F0558",
000673 => x"EBFFFE75",
000674 => x"EAFFFF6D",
000675 => x"E1A00004",
000676 => x"EBFFFD9F",
000677 => x"E59F0548",
000678 => x"EBFFFE70",
000679 => x"E59F0544",
000680 => x"EBFFFE6E",
000681 => x"EAFFFF66",
000682 => x"E5DD3011",
000683 => x"E3530042",
000684 => x"1AFFFF91",
000685 => x"E3500052",
000686 => x"1AFFFF8F",
000687 => x"E1A01004",
000688 => x"E3A02004",
000689 => x"E2433040",
000690 => x"E2800020",
000691 => x"E58D5000",
000692 => x"EBFFFDCB",
000693 => x"E1A01004",
000694 => x"E5CD000F",
000695 => x"E3A02005",
000696 => x"E3A03002",
000697 => x"E3A00072",
000698 => x"E58D5000",
000699 => x"EBFFFDC4",
000700 => x"E1A01004",
000701 => x"E5CD0010",
000702 => x"E3A02006",
000703 => x"E3A03002",
000704 => x"E3A00072",
000705 => x"E58D5000",
000706 => x"EBFFFDBD",
000707 => x"E1A01004",
000708 => x"E5CD0011",
000709 => x"E3A02007",
000710 => x"E3A03002",
000711 => x"E3A00072",
000712 => x"E58D5000",
000713 => x"EBFFFDB6",
000714 => x"E5CD0012",
000715 => x"E1A0000A",
000716 => x"EBFFFF0A",
000717 => x"E3700004",
000718 => x"E58D0014",
000719 => x"0A000024",
000720 => x"E1A06005",
000721 => x"E2852008",
000722 => x"E1A01004",
000723 => x"E3A03002",
000724 => x"E3A00072",
000725 => x"E58D6000",
000726 => x"EBFFFDA9",
000727 => x"E2852009",
000728 => x"E5CD000F",
000729 => x"E1A01004",
000730 => x"E3A03002",
000731 => x"E3A00072",
000732 => x"E58D6000",
000733 => x"EBFFFDA2",
000734 => x"E285200A",
000735 => x"E5CD0010",
000736 => x"E1A01004",
000737 => x"E3A03002",
000738 => x"E3A00072",
000739 => x"E58D6000",
000740 => x"EBFFFD9B",
000741 => x"E285200B",
000742 => x"E3A03002",
000743 => x"E5CD0011",
000744 => x"E1A01004",
000745 => x"E3A00072",
000746 => x"E58D6000",
000747 => x"EBFFFD94",
000748 => x"E5CD0012",
000749 => x"E1A0000A",
000750 => x"EBFFFEE8",
000751 => x"E4850004",
000752 => x"E59D3014",
000753 => x"E2833004",
000754 => x"E1530005",
000755 => x"13550902",
000756 => x"3AFFFFDB",
000757 => x"E59F0410",
000758 => x"EBFFFE20",
000759 => x"EAFFFF4A",
000760 => x"E3740001",
000761 => x"0AFFFF16",
000762 => x"E3540030",
000763 => x"0A000004",
000764 => x"E20400FF",
000765 => x"EBFFFD46",
000766 => x"E59F03F0",
000767 => x"EBFFFE17",
000768 => x"EAFFFF0F",
000769 => x"E1A00004",
000770 => x"EBFFFD41",
000771 => x"EAFFFF3E",
000772 => x"E1A00004",
000773 => x"EBFFFD3E",
000774 => x"E59F03D4",
000775 => x"EBFFFE0F",
000776 => x"EBFFFD35",
000777 => x"E3700001",
000778 => x"0AFFFFFC",
000779 => x"EBFFFD32",
000780 => x"E3700001",
000781 => x"1AFFFFFC",
000782 => x"E3A05301",
000783 => x"E5950000",
000784 => x"E1A01009",
000785 => x"E3A02008",
000786 => x"EBFFFE32",
000787 => x"E5DD0006",
000788 => x"E3500000",
000789 => x"0A000005",
000790 => x"E3A04000",
000791 => x"E2844001",
000792 => x"EBFFFD2B",
000793 => x"E7D40009",
000794 => x"E3500000",
000795 => x"1AFFFFFA",
000796 => x"E3A00020",
000797 => x"EBFFFD26",
000798 => x"EBFFFD1F",
000799 => x"E3700001",
000800 => x"1A000005",
000801 => x"E3A03301",
000802 => x"E2833E9E",
000803 => x"E2855004",
000804 => x"E2833004",
000805 => x"E1550003",
000806 => x"1AFFFFE7",
000807 => x"E59F0354",
000808 => x"EBFFFDEE",
000809 => x"EAFFFEE6",
000810 => x"E3540035",
000811 => x"0A000087",
000812 => x"E3540061",
000813 => x"1AFFFFCD",
000814 => x"E1A00004",
000815 => x"EBFFFD14",
000816 => x"E59F0334",
000817 => x"EBFFFDE5",
000818 => x"E59F0330",
000819 => x"EBFFFDE3",
000820 => x"E59F032C",
000821 => x"EBFFFDE1",
000822 => x"EAFFFED9",
000823 => x"E59F0324",
000824 => x"EBFFFDDE",
000825 => x"E1A0000A",
000826 => x"E3A01004",
000827 => x"E3A02000",
000828 => x"EBFFFDE8",
000829 => x"E5DD300F",
000830 => x"E3530053",
000831 => x"1A000002",
000832 => x"E5DD2010",
000833 => x"E352004D",
000834 => x"0A000004",
000835 => x"E59F02F8",
000836 => x"EBFFFDD2",
000837 => x"E59F02F4",
000838 => x"EBFFFDD0",
000839 => x"EAFFFEC8",
000840 => x"E5DD1011",
000841 => x"E3510042",
000842 => x"1AFFFFF7",
000843 => x"E5DD0012",
000844 => x"E3500052",
000845 => x"1AFFFFF4",
000846 => x"E3A04000",
000847 => x"E5C43000",
000848 => x"E1A00000",
000849 => x"E5C42001",
000850 => x"E1A00000",
000851 => x"E5C41002",
000852 => x"E1A00000",
000853 => x"E5C40003",
000854 => x"E1A00000",
000855 => x"E241103E",
000856 => x"E1A0000A",
000857 => x"E1A02004",
000858 => x"EBFFFDCA",
000859 => x"E5DD300F",
000860 => x"E5C43004",
000861 => x"E5DD2010",
000862 => x"E5C42005",
000863 => x"E5DD3011",
000864 => x"E5C43006",
000865 => x"E5DD2012",
000866 => x"E1A0000A",
000867 => x"E5C42007",
000868 => x"EBFFFE72",
000869 => x"E3A03CFF",
000870 => x"E28330FC",
000871 => x"E1500003",
000872 => x"E1A05000",
000873 => x"8A000076",
000874 => x"E3700004",
000875 => x"12844008",
000876 => x"1280600B",
000877 => x"0A000006",
000878 => x"EBFFFCCF",
000879 => x"E3700001",
000880 => x"0AFFFFFC",
000881 => x"E1560004",
000882 => x"E5C40000",
000883 => x"E2844001",
000884 => x"1AFFFFF8",
000885 => x"E59F0238",
000886 => x"EBFFFDA0",
000887 => x"E59F0234",
000888 => x"EBFFFD9E",
000889 => x"E375000C",
000890 => x"0A00000F",
000891 => x"E3A04000",
000892 => x"E285700C",
000893 => x"E1A06004",
000894 => x"E5D45000",
000895 => x"E3A00077",
000896 => x"E1A01008",
000897 => x"E1A02006",
000898 => x"E3A03002",
000899 => x"E58D5000",
000900 => x"EBFFFCFB",
000901 => x"E3500000",
000902 => x"1AFFFFF7",
000903 => x"E2844001",
000904 => x"E1540007",
000905 => x"E1A06004",
000906 => x"1AFFFFF2",
000907 => x"E59F01E8",
000908 => x"EBFFFD8A",
000909 => x"EAFFFFB6",
000910 => x"E1A00004",
000911 => x"EBFFFCB4",
000912 => x"EBFFFE17",
000913 => x"EAFFFE7E",
000914 => x"E5DD3011",
000915 => x"E3530042",
000916 => x"1AFFFF0A",
000917 => x"E5DD3012",
000918 => x"E3530052",
000919 => x"1AFFFF07",
000920 => x"E3A01004",
000921 => x"E3A02000",
000922 => x"E1A0000A",
000923 => x"EBFFFD89",
000924 => x"E1A0000A",
000925 => x"EBFFFE39",
000926 => x"E3700008",
000927 => x"E58D0014",
000928 => x"8A00003C",
000929 => x"E2804301",
000930 => x"E2844004",
000931 => x"E3540301",
000932 => x"0A000009",
000933 => x"E3A05301",
000934 => x"E3A01004",
000935 => x"E3A02000",
000936 => x"E1A0000A",
000937 => x"EBFFFD7B",
000938 => x"E1A0000A",
000939 => x"EBFFFE2B",
000940 => x"E4850004",
000941 => x"E1550004",
000942 => x"1AFFFFF6",
000943 => x"E59F015C",
000944 => x"EBFFFD66",
000945 => x"E59F0158",
000946 => x"EBFFFD64",
000947 => x"EAFFFE5C",
000948 => x"E1A00004",
000949 => x"EBFFFC8E",
000950 => x"E59F0148",
000951 => x"EBFFFD5F",
000952 => x"E1A0000A",
000953 => x"E3A01002",
000954 => x"E3A02001",
000955 => x"EBFFFD69",
000956 => x"E1A0000A",
000957 => x"E3A01002",
000958 => x"EBFFFDCE",
000959 => x"E21060FF",
000960 => x"0AFFFEAD",
000961 => x"E59F0120",
000962 => x"EBFFFD54",
000963 => x"E59F011C",
000964 => x"EBFFFD52",
000965 => x"EBFFFC78",
000966 => x"E3700001",
000967 => x"0AFFFFFC",
000968 => x"EBFFFC75",
000969 => x"E3700001",
000970 => x"1AFFFFFC",
000971 => x"E3A05000",
000972 => x"EA000001",
000973 => x"E3540000",
000974 => x"AA000014",
000975 => x"E3A0C000",
000976 => x"E1A02005",
000977 => x"E1A01006",
000978 => x"E3A03002",
000979 => x"E3A00072",
000980 => x"E58DC000",
000981 => x"EBFFFCAA",
000982 => x"E1A04000",
000983 => x"EBFFFC66",
000984 => x"E3700001",
000985 => x"E1A00004",
000986 => x"0AFFFFF1",
000987 => x"E59F00C0",
000988 => x"EBFFFD3A",
000989 => x"EAFFFF48",
000990 => x"E59F00B8",
000991 => x"EBFFFD37",
000992 => x"EAFFFE2F",
000993 => x"E59F00B0",
000994 => x"EBFFFD34",
000995 => x"EAFFFE2C",
000996 => x"EBFFFC5F",
000997 => x"E3A03801",
000998 => x"E2855001",
000999 => x"E2433001",
001000 => x"E1550003",
001001 => x"1AFFFFE4",
001002 => x"EAFFFF3B",
001003 => x"000114B8",
001004 => x"000114D0",
001005 => x"000114D8",
001006 => x"00011694",
001007 => x"000116F8",
001008 => x"00011A58",
001009 => x"00011A7C",
001010 => x"00011AAC",
001011 => x"00011AD0",
001012 => x"00011638",
001013 => x"00011674",
001014 => x"00011724",
001015 => x"000114E8",
001016 => x"000115A4",
001017 => x"000119DC",
001018 => x"00011A0C",
001019 => x"000116E4",
001020 => x"00011A34",
001021 => x"000115CC",
001022 => x"00011614",
001023 => x"000118F8",
001024 => x"0001192C",
001025 => x"00011998",
001026 => x"00011744",
001027 => x"00011810",
001028 => x"00011A28",
001029 => x"000117C8",
001030 => x"000117E0",
001031 => x"00011800",
001032 => x"00011584",
001033 => x"00011594",
001034 => x"00011834",
001035 => x"00011870",
001036 => x"000118B0",
001037 => x"00011AEC",
001038 => x"0001155C",
001039 => x"000117A4",
001040 => x"E10F3000",
001041 => x"E3C330C0",
001042 => x"E129F003",
001043 => x"E1A0F00E",
001044 => x"E10F3000",
001045 => x"E38330C0",
001046 => x"E129F003",
001047 => x"E1A0F00E",
001048 => x"00000000",
001049 => x"0D0A0D0A",
001050 => x"0D0A2B2D",
001051 => x"2D2D2D2D",
001052 => x"2D2D2D2D",
001053 => x"2D2D2D2D",
001054 => x"2D2D2D2D",
001055 => x"2D2D2D2D",
001056 => x"2D2D2D2D",
001057 => x"2D2D2D2D",
001058 => x"2D2D2D2D",
001059 => x"2D2D2D2D",
001060 => x"2D2D2D2D",
001061 => x"2D2D2D2D",
001062 => x"2D2D2D2D",
001063 => x"2D2D2D2D",
001064 => x"2D2D2D2D",
001065 => x"2D2D2D2D",
001066 => x"2D2D2D2B",
001067 => x"0D0A0000",
001068 => x"7C202020",
001069 => x"203C3C3C",
001070 => x"2053544F",
001071 => x"524D2043",
001072 => x"6F726520",
001073 => x"50726F63",
001074 => x"6573736F",
001075 => x"72205379",
001076 => x"7374656D",
001077 => x"202D2042",
001078 => x"79205374",
001079 => x"65706861",
001080 => x"6E204E6F",
001081 => x"6C74696E",
001082 => x"67203E3E",
001083 => x"3E202020",
001084 => x"207C0D0A",
001085 => x"00000000",
001086 => x"2B2D2D2D",
001087 => x"2D2D2D2D",
001088 => x"2D2D2D2D",
001089 => x"2D2D2D2D",
001090 => x"2D2D2D2D",
001091 => x"2D2D2D2D",
001092 => x"2D2D2D2D",
001093 => x"2D2D2D2D",
001094 => x"2D2D2D2D",
001095 => x"2D2D2D2D",
001096 => x"2D2D2D2D",
001097 => x"2D2D2D2D",
001098 => x"2D2D2D2D",
001099 => x"2D2D2D2D",
001100 => x"2D2D2D2D",
001101 => x"2D2D2D2D",
001102 => x"2D2B0D0A",
001103 => x"00000000",
001104 => x"7C202020",
001105 => x"20202020",
001106 => x"2020426F",
001107 => x"6F746C6F",
001108 => x"61646572",
001109 => x"20666F72",
001110 => x"2053544F",
001111 => x"524D2053",
001112 => x"6F432020",
001113 => x"20566572",
001114 => x"73696F6E",
001115 => x"3A203230",
001116 => x"31323035",
001117 => x"32342D44",
001118 => x"20202020",
001119 => x"20202020",
001120 => x"207C0D0A",
001121 => x"00000000",
001122 => x"7C202020",
001123 => x"20202020",
001124 => x"20202020",
001125 => x"20202020",
001126 => x"436F6E74",
001127 => x"6163743A",
001128 => x"2073746E",
001129 => x"6F6C7469",
001130 => x"6E674067",
001131 => x"6F6F676C",
001132 => x"656D6169",
001133 => x"6C2E636F",
001134 => x"6D202020",
001135 => x"20202020",
001136 => x"20202020",
001137 => x"20202020",
001138 => x"207C0D0A",
001139 => x"00000000",
001140 => x"2B2D2D2D",
001141 => x"2D2D2D2D",
001142 => x"2D2D2D2D",
001143 => x"2D2D2D2D",
001144 => x"2D2D2D2D",
001145 => x"2D2D2D2D",
001146 => x"2D2D2D2D",
001147 => x"2D2D2D2D",
001148 => x"2D2D2D2D",
001149 => x"2D2D2D2D",
001150 => x"2D2D2D2D",
001151 => x"2D2D2D2D",
001152 => x"2D2D2D2D",
001153 => x"2D2D2D2D",
001154 => x"2D2D2D2D",
001155 => x"2D2D2D2D",
001156 => x"2D2B0D0A",
001157 => x"0D0A0000",
001158 => x"636F6E6E",
001159 => x"65637465",
001160 => x"6420746F",
001161 => x"20493243",
001162 => x"5F434F4E",
001163 => x"54524F4C",
001164 => x"4C45525F",
001165 => x"302C206F",
001166 => x"70657261",
001167 => x"74696E67",
001168 => x"20667265",
001169 => x"7175656E",
001170 => x"63792069",
001171 => x"73203130",
001172 => x"306B487A",
001173 => x"2C0D0A00",
001174 => x"6D617869",
001175 => x"6D756D20",
001176 => x"45455052",
001177 => x"4F4D2073",
001178 => x"697A6520",
001179 => x"3D203635",
001180 => x"35333620",
001181 => x"62797465",
001182 => x"203D3E20",
001183 => x"31362062",
001184 => x"69742061",
001185 => x"64647265",
001186 => x"73736573",
001187 => x"2C0D0A00",
001188 => x"66697865",
001189 => x"6420626F",
001190 => x"6F742064",
001191 => x"65766963",
001192 => x"65206164",
001193 => x"64726573",
001194 => x"733A2030",
001195 => x"7841300D",
001196 => x"0A0D0A00",
001197 => x"426F6F74",
001198 => x"20454550",
001199 => x"524F4D3A",
001200 => x"20323478",
001201 => x"786E6E6E",
001202 => x"20286C69",
001203 => x"6B652032",
001204 => x"34414136",
001205 => x"34292C20",
001206 => x"37206269",
001207 => x"74206164",
001208 => x"64726573",
001209 => x"73202B20",
001210 => x"646F6E74",
001211 => x"2D636172",
001212 => x"65206269",
001213 => x"742C0D0A",
001214 => x"00000000",
001215 => x"203C2057",
001216 => x"656C636F",
001217 => x"6D652074",
001218 => x"6F207468",
001219 => x"65205354",
001220 => x"4F524D20",
001221 => x"536F4320",
001222 => x"626F6F74",
001223 => x"6C6F6164",
001224 => x"65722063",
001225 => x"6F6E736F",
001226 => x"6C652120",
001227 => x"3E0D0A20",
001228 => x"3C205365",
001229 => x"6C656374",
001230 => x"20616E20",
001231 => x"6F706572",
001232 => x"6174696F",
001233 => x"6E206672",
001234 => x"6F6D2074",
001235 => x"6865206D",
001236 => x"656E7520",
001237 => x"62656C6F",
001238 => x"77206F72",
001239 => x"20707265",
001240 => x"7373203E",
001241 => x"0D0A0000",
001242 => x"203C2074",
001243 => x"68652062",
001244 => x"6F6F7420",
001245 => x"6B657920",
001246 => x"666F7220",
001247 => x"696D6D65",
001248 => x"64696174",
001249 => x"65206170",
001250 => x"706C6963",
001251 => x"6174696F",
001252 => x"6E207374",
001253 => x"6172742E",
001254 => x"203E0D0A",
001255 => x"0D0A0000",
001256 => x"2030202D",
001257 => x"20626F6F",
001258 => x"74206672",
001259 => x"6F6D2063",
001260 => x"6F726520",
001261 => x"52414D20",
001262 => x"28737461",
001263 => x"72742061",
001264 => x"70706C69",
001265 => x"63617469",
001266 => x"6F6E290D",
001267 => x"0A203120",
001268 => x"2D207072",
001269 => x"6F677261",
001270 => x"6D20636F",
001271 => x"72652052",
001272 => x"414D2076",
001273 => x"69612055",
001274 => x"4152545F",
001275 => x"300D0A20",
001276 => x"32202D20",
001277 => x"636F7265",
001278 => x"2052414D",
001279 => x"2064756D",
001280 => x"700D0A00",
001281 => x"2033202D",
001282 => x"20626F6F",
001283 => x"74206672",
001284 => x"6F6D2049",
001285 => x"32432045",
001286 => x"4550524F",
001287 => x"4D0D0A20",
001288 => x"34202D20",
001289 => x"70726F67",
001290 => x"72616D20",
001291 => x"49324320",
001292 => x"45455052",
001293 => x"4F4D2076",
001294 => x"69612055",
001295 => x"4152545F",
001296 => x"300D0A20",
001297 => x"35202D20",
001298 => x"73686F77",
001299 => x"20636F6E",
001300 => x"74656E74",
001301 => x"206F6620",
001302 => x"49324320",
001303 => x"45455052",
001304 => x"4F4D0D0A",
001305 => x"00000000",
001306 => x"2061202D",
001307 => x"20617574",
001308 => x"6F6D6174",
001309 => x"69632062",
001310 => x"6F6F7420",
001311 => x"636F6E66",
001312 => x"69677572",
001313 => x"6174696F",
001314 => x"6E0D0A20",
001315 => x"68202D20",
001316 => x"68656C70",
001317 => x"0D0A2072",
001318 => x"202D2072",
001319 => x"65737461",
001320 => x"72742073",
001321 => x"79737465",
001322 => x"6D0D0A0D",
001323 => x"0A53656C",
001324 => x"6563743A",
001325 => x"20000000",
001326 => x"41646472",
001327 => x"65737320",
001328 => x"6F662061",
001329 => x"64725F62",
001330 => x"75666665",
001331 => x"723A2000",
001332 => x"200A0D20",
001333 => x"00000000",
001334 => x"204C6F61",
001335 => x"64204164",
001336 => x"64726573",
001337 => x"733A2000",
001338 => x"0D0A0D0A",
001339 => x"4170706C",
001340 => x"69636174",
001341 => x"696F6E20",
001342 => x"77696C6C",
001343 => x"20737461",
001344 => x"72742061",
001345 => x"75746F6D",
001346 => x"61746963",
001347 => x"616C6C79",
001348 => x"20616674",
001349 => x"65722064",
001350 => x"6F776E6C",
001351 => x"6F61642E",
001352 => x"0D0A2D3E",
001353 => x"20576169",
001354 => x"74696E67",
001355 => x"20666F72",
001356 => x"20277374",
001357 => x"6F726D5F",
001358 => x"70726F67",
001359 => x"72616D2E",
001360 => x"62696E27",
001361 => x"20696E20",
001362 => x"62797465",
001363 => x"2D737472",
001364 => x"65616D20",
001365 => x"6D6F6465",
001366 => x"2E2E2E00",
001367 => x"20534452",
001368 => x"414D2045",
001369 => x"52524F52",
001370 => x"21205072",
001371 => x"6F677261",
001372 => x"6D206669",
001373 => x"6C652074",
001374 => x"6F6F2062",
001375 => x"6967210D",
001376 => x"0A0D0A00",
001377 => x"446F6E65",
001378 => x"204C6F61",
001379 => x"64696E67",
001380 => x"210D0A00",
001381 => x"4C415354",
001382 => x"20414444",
001383 => x"52455353",
001384 => x"3A000000",
001385 => x"20496E76",
001386 => x"616C6964",
001387 => x"2070726F",
001388 => x"6772616D",
001389 => x"6D696E67",
001390 => x"2066696C",
001391 => x"65210D0A",
001392 => x"0D0A5365",
001393 => x"6C656374",
001394 => x"3A200000",
001395 => x"0D0A0D0A",
001396 => x"41626F72",
001397 => x"74206475",
001398 => x"6D70696E",
001399 => x"67206279",
001400 => x"20707265",
001401 => x"7373696E",
001402 => x"6720616E",
001403 => x"79206B65",
001404 => x"792E0D0A",
001405 => x"50726573",
001406 => x"7320616E",
001407 => x"79206B65",
001408 => x"7920746F",
001409 => x"20636F6E",
001410 => x"74696E75",
001411 => x"652E0D0A",
001412 => x"0D0A0000",
001413 => x"0D0A0D0A",
001414 => x"44756D70",
001415 => x"696E6720",
001416 => x"636F6D70",
001417 => x"6C657465",
001418 => x"642E0D0A",
001419 => x"0D0A5365",
001420 => x"6C656374",
001421 => x"3A200000",
001422 => x"0D0A0D0A",
001423 => x"456E7465",
001424 => x"72206465",
001425 => x"76696365",
001426 => x"20616464",
001427 => x"72657373",
001428 => x"20283278",
001429 => x"20686578",
001430 => x"5F636861",
001431 => x"72732C20",
001432 => x"73657420",
001433 => x"4C534220",
001434 => x"746F2027",
001435 => x"3027293A",
001436 => x"20000000",
001437 => x"20496E76",
001438 => x"616C6964",
001439 => x"20616464",
001440 => x"72657373",
001441 => x"210D0A0D",
001442 => x"0A53656C",
001443 => x"6563743A",
001444 => x"20000000",
001445 => x"0D0A4170",
001446 => x"706C6963",
001447 => x"6174696F",
001448 => x"6E207769",
001449 => x"6C6C2073",
001450 => x"74617274",
001451 => x"20617574",
001452 => x"6F6D6174",
001453 => x"6963616C",
001454 => x"6C792061",
001455 => x"66746572",
001456 => x"2075706C",
001457 => x"6F61642E",
001458 => x"0D0A2D3E",
001459 => x"204C6F61",
001460 => x"64696E67",
001461 => x"20626F6F",
001462 => x"7420696D",
001463 => x"6167652E",
001464 => x"2E2E0000",
001465 => x"2055706C",
001466 => x"6F616420",
001467 => x"636F6D70",
001468 => x"6C657465",
001469 => x"0D0A0000",
001470 => x"20496E76",
001471 => x"616C6964",
001472 => x"20626F6F",
001473 => x"74206465",
001474 => x"76696365",
001475 => x"206F7220",
001476 => x"66696C65",
001477 => x"210D0A0D",
001478 => x"0A53656C",
001479 => x"6563743A",
001480 => x"20000000",
001481 => x"0D0A496E",
001482 => x"76616C69",
001483 => x"64206164",
001484 => x"64726573",
001485 => x"73210D0A",
001486 => x"0D0A5365",
001487 => x"6C656374",
001488 => x"3A200000",
001489 => x"0D0A4461",
001490 => x"74612077",
001491 => x"696C6C20",
001492 => x"6F766572",
001493 => x"77726974",
001494 => x"65205241",
001495 => x"4D20636F",
001496 => x"6E74656E",
001497 => x"74210D0A",
001498 => x"2D3E2057",
001499 => x"61697469",
001500 => x"6E672066",
001501 => x"6F722027",
001502 => x"73746F72",
001503 => x"6D5F7072",
001504 => x"6F677261",
001505 => x"6D2E6269",
001506 => x"6E272069",
001507 => x"6E206279",
001508 => x"74652D73",
001509 => x"74726561",
001510 => x"6D206D6F",
001511 => x"64652E2E",
001512 => x"2E000000",
001513 => x"20455252",
001514 => x"4F522120",
001515 => x"50726F67",
001516 => x"72616D20",
001517 => x"66696C65",
001518 => x"20746F6F",
001519 => x"20626967",
001520 => x"210D0A0D",
001521 => x"0A000000",
001522 => x"20446F77",
001523 => x"6E6C6F61",
001524 => x"6420636F",
001525 => x"6D706C65",
001526 => x"7465640D",
001527 => x"0A000000",
001528 => x"57726974",
001529 => x"696E6720",
001530 => x"62756666",
001531 => x"65722074",
001532 => x"6F206932",
001533 => x"63204545",
001534 => x"50524F4D",
001535 => x"2E2E2E00",
001536 => x"20436F6D",
001537 => x"706C6574",
001538 => x"65640D0A",
001539 => x"0D0A0000",
001540 => x"20496E76",
001541 => x"616C6964",
001542 => x"20626F6F",
001543 => x"74206465",
001544 => x"76696365",
001545 => x"206F7220",
001546 => x"66696C65",
001547 => x"210D0A0D",
001548 => x"0A000000",
001549 => x"0D0A0D0A",
001550 => x"456E7465",
001551 => x"72206465",
001552 => x"76696365",
001553 => x"20616464",
001554 => x"72657373",
001555 => x"20283220",
001556 => x"6865782D",
001557 => x"63686172",
001558 => x"732C2073",
001559 => x"6574204C",
001560 => x"53422074",
001561 => x"6F202730",
001562 => x"27293A20",
001563 => x"00000000",
001564 => x"0D0A0D0A",
001565 => x"41626F72",
001566 => x"74206475",
001567 => x"6D70696E",
001568 => x"67206279",
001569 => x"20707265",
001570 => x"7373696E",
001571 => x"6720616E",
001572 => x"79206B65",
001573 => x"792E2049",
001574 => x"66206E6F",
001575 => x"20646174",
001576 => x"61206973",
001577 => x"2073686F",
001578 => x"776E2C0D",
001579 => x"0A000000",
001580 => x"74686520",
001581 => x"73656C65",
001582 => x"63746564",
001583 => x"20646576",
001584 => x"69636520",
001585 => x"6973206E",
001586 => x"6F742072",
001587 => x"6573706F",
001588 => x"6E64696E",
001589 => x"672E2050",
001590 => x"72657373",
001591 => x"20616E79",
001592 => x"206B6579",
001593 => x"20746F20",
001594 => x"636F6E74",
001595 => x"696E7565",
001596 => x"2E0D0A0D",
001597 => x"0A000000",
001598 => x"0D0A0D0A",
001599 => x"4175746F",
001600 => x"6D617469",
001601 => x"6320626F",
001602 => x"6F742063",
001603 => x"6F6E6669",
001604 => x"67757261",
001605 => x"74696F6E",
001606 => x"20666F72",
001607 => x"20706F77",
001608 => x"65722D75",
001609 => x"703A0D0A",
001610 => x"00000000",
001611 => x"5B333231",
001612 => x"305D2063",
001613 => x"6F6E6669",
001614 => x"67757261",
001615 => x"74696F6E",
001616 => x"20444950",
001617 => x"20737769",
001618 => x"7463680D",
001619 => x"0A203030",
001620 => x"3030202D",
001621 => x"20537461",
001622 => x"72742062",
001623 => x"6F6F746C",
001624 => x"6F616465",
001625 => x"7220636F",
001626 => x"6E736F6C",
001627 => x"650D0A20",
001628 => x"30303031",
001629 => x"202D2041",
001630 => x"75746F6D",
001631 => x"61746963",
001632 => x"20626F6F",
001633 => x"74206672",
001634 => x"6F6D2063",
001635 => x"6F726520",
001636 => x"52414D0D",
001637 => x"0A000000",
001638 => x"20303031",
001639 => x"30202D20",
001640 => x"4175746F",
001641 => x"6D617469",
001642 => x"6320626F",
001643 => x"6F742066",
001644 => x"726F6D20",
001645 => x"49324320",
001646 => x"45455052",
001647 => x"4F4D2028",
001648 => x"41646472",
001649 => x"65737320",
001650 => x"30784130",
001651 => x"290D0A0D",
001652 => x"0A53656C",
001653 => x"6563743A",
001654 => x"20000000",
001655 => x"0D0A0D0A",
001656 => x"5765276C",
001657 => x"6C207365",
001658 => x"6E642079",
001659 => x"6F752062",
001660 => x"61636B20",
001661 => x"2D20746F",
001662 => x"20746865",
001663 => x"20667574",
001664 => x"75726521",
001665 => x"2E0D0A0D",
001666 => x"0A000000",
001667 => x"202D2044",
001668 => x"6F63746F",
001669 => x"7220456D",
001670 => x"6D657420",
001671 => x"4C2E2042",
001672 => x"726F776E",
001673 => x"0D0A0D0A",
001674 => x"53656C65",
001675 => x"63743A20",
001676 => x"00000000",
001677 => x"20496E76",
001678 => x"616C6964",
001679 => x"206F7065",
001680 => x"72617469",
001681 => x"6F6E210D",
001682 => x"0A547279",
001683 => x"20616761",
001684 => x"696E3A20",
001685 => x"00000000",
001686 => x"0D0A0D0A",
001687 => x"2D3E2053",
001688 => x"74617274",
001689 => x"696E6720",
001690 => x"6170706C",
001691 => x"69636174",
001692 => x"696F6E2E",
001693 => x"2E2E0D0A",
001694 => x"0D0A0000",
001695 => x"0D0A0D0A",
001696 => x"2D3E2064",
001697 => x"69736162",
001698 => x"6C652077",
001699 => x"72697465",
001700 => x"2D746872",
001701 => x"6F756768",
001702 => x"20737472",
001703 => x"61746567",
001704 => x"792E2E2E",
001705 => x"0D0A0D0A",
001706 => x"00000000",
001707 => x"0D0A0D0A",
001708 => x"2D3E206A",
001709 => x"756D7020",
001710 => x"746F2061",
001711 => x"70706C69",
001712 => x"63617469",
001713 => x"6F6E2E2E",
001714 => x"2E0D0A0D",
001715 => x"0A000000",
001716 => x"21217368",
001717 => x"6F756C64",
001718 => x"206E6F74",
001719 => x"20626520",
001720 => x"68657265",
001721 => x"21210D0A",
001722 => x"00000000",
001723 => x"0D0A0D0A",
001724 => x"41626F72",
001725 => x"74656421",
001726 => x"00000000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;