-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
000000 => x"EA000006",
000001 => x"EAFFFFFE",
000002 => x"EAFFFFFE",
000003 => x"EAFFFFFE",
000004 => x"EAFFFFFE",
000005 => x"E1A00000",
000006 => x"EAFFFFFE",
000007 => x"EAFFFFFE",
000008 => x"E59F0034",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA00C",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"EAFFFFFE",
000023 => x"00002000",
000024 => x"00010778",
000025 => x"E3E03A0F",
000026 => x"E5131FFB",
000027 => x"E20020FF",
000028 => x"E3A00001",
000029 => x"E0010210",
000030 => x"E1A0F00E",
000031 => x"E3E03A0F",
000032 => x"E5130FFB",
000033 => x"E1A0F00E",
000034 => x"E3E01A0F",
000035 => x"E5113FFF",
000036 => x"E20000FF",
000037 => x"E3A02001",
000038 => x"E1833012",
000039 => x"E5013FFF",
000040 => x"E1A0F00E",
000041 => x"E20000FF",
000042 => x"E3A02001",
000043 => x"E1A02012",
000044 => x"E3E01A0F",
000045 => x"E5113FFF",
000046 => x"E1E02002",
000047 => x"E0033002",
000048 => x"E5013FFF",
000049 => x"E1A0F00E",
000050 => x"E3E01A0F",
000051 => x"E5113FFF",
000052 => x"E20000FF",
000053 => x"E3A02001",
000054 => x"E0233012",
000055 => x"E5013FFF",
000056 => x"E1A0F00E",
000057 => x"E3E03A0F",
000058 => x"E5030FFF",
000059 => x"E1A0F00E",
000060 => x"E20000FF",
000061 => x"E3500007",
000062 => x"E92D4010",
000063 => x"E3A0C000",
000064 => x"E3E0E0FF",
000065 => x"E20110FF",
000066 => x"8A000011",
000067 => x"E2403004",
000068 => x"E20330FF",
000069 => x"E3500003",
000070 => x"E1A0E183",
000071 => x"E3E04A0F",
000072 => x"E1A0C180",
000073 => x"9A000007",
000074 => x"E3A030FF",
000075 => x"E1A03E13",
000076 => x"E5142F8B",
000077 => x"E1E03003",
000078 => x"E0022003",
000079 => x"E1822E11",
000080 => x"E5042F8B",
000081 => x"E8BD8010",
000082 => x"E3A030FF",
000083 => x"E1A03C13",
000084 => x"E1E0E003",
000085 => x"E3E02A0F",
000086 => x"E5123F8F",
000087 => x"E003300E",
000088 => x"E1833C11",
000089 => x"E5023F8F",
000090 => x"E8BD8010",
000091 => x"E20000FF",
000092 => x"E3500007",
000093 => x"E3A02000",
000094 => x"8A00000A",
000095 => x"E2403004",
000096 => x"E3500003",
000097 => x"E20320FF",
000098 => x"9A000005",
000099 => x"E3E03A0F",
000100 => x"E5130F8B",
000101 => x"E1A02182",
000102 => x"E1A00230",
000103 => x"E20000FF",
000104 => x"E1A0F00E",
000105 => x"E1A02180",
000106 => x"E3E03A0F",
000107 => x"E5130F8F",
000108 => x"E1A00230",
000109 => x"E20000FF",
000110 => x"E1A0F00E",
000111 => x"E3E02A0F",
000112 => x"E5123FE3",
000113 => x"E3130002",
000114 => x"E3E00000",
000115 => x"15120FE7",
000116 => x"E1A0F00E",
000117 => x"E3E02A0F",
000118 => x"E5123FE3",
000119 => x"E3130001",
000120 => x"0AFFFFFC",
000121 => x"E20030FF",
000122 => x"E5023FE7",
000123 => x"E1A0F00E",
000124 => x"E20000FF",
000125 => x"E3500001",
000126 => x"E3812B01",
000127 => x"03E03A0F",
000128 => x"E3811B09",
000129 => x"13E03A0F",
000130 => x"05031FCF",
000131 => x"15032FCF",
000132 => x"E1A0F00E",
000133 => x"E3E03A0F",
000134 => x"E5030FCB",
000135 => x"E1A0F00E",
000136 => x"E3E02A0F",
000137 => x"E5123FCF",
000138 => x"E3130C01",
000139 => x"1AFFFFFC",
000140 => x"E5020FBF",
000141 => x"E5123FCF",
000142 => x"E3833C01",
000143 => x"E5023FCF",
000144 => x"E3E02A0F",
000145 => x"E5123FCF",
000146 => x"E3130C01",
000147 => x"1AFFFFFC",
000148 => x"E5120FBF",
000149 => x"E1A0F00E",
000150 => x"E3E01A0F",
000151 => x"E5113FC7",
000152 => x"E20000FF",
000153 => x"E3A02001",
000154 => x"E1833012",
000155 => x"E5013FC7",
000156 => x"E1A0F00E",
000157 => x"E20000FF",
000158 => x"E3A02001",
000159 => x"E1A02012",
000160 => x"E3E01A0F",
000161 => x"E5113FC7",
000162 => x"E1E02002",
000163 => x"E0033002",
000164 => x"E5013FC7",
000165 => x"E1A0F00E",
000166 => x"E3E02A0F",
000167 => x"E5123F97",
000168 => x"E1A01420",
000169 => x"E3C33080",
000170 => x"E5023F97",
000171 => x"E5020F9F",
000172 => x"E5021F9B",
000173 => x"E5123F97",
000174 => x"E3833080",
000175 => x"E5023F97",
000176 => x"E1A0F00E",
000177 => x"E92D4030",
000178 => x"E3A0C090",
000179 => x"E20140FE",
000180 => x"E3E0EA0F",
000181 => x"E5DD500F",
000182 => x"E20000FF",
000183 => x"E50E4F93",
000184 => x"E20110FF",
000185 => x"E50ECFAF",
000186 => x"E1A04002",
000187 => x"E203C0FF",
000188 => x"E51E3FAF",
000189 => x"E3130002",
000190 => x"1AFFFFFC",
000191 => x"E51E3FAF",
000192 => x"E3130080",
000193 => x"13E00000",
000194 => x"18BD8030",
000195 => x"E35C0000",
000196 => x"0A000012",
000197 => x"E24C3001",
000198 => x"E203C0FF",
000199 => x"E35C0001",
000200 => x"01A02424",
000201 => x"03E03A0F",
000202 => x"13E03A0F",
000203 => x"05032F93",
000204 => x"15034F93",
000205 => x"E3E02A0F",
000206 => x"E3A03010",
000207 => x"E5023FAF",
000208 => x"E5123FAF",
000209 => x"E3130002",
000210 => x"1AFFFFFC",
000211 => x"E5123FAF",
000212 => x"E3130080",
000213 => x"0AFFFFEC",
000214 => x"E3E00001",
000215 => x"E8BD8030",
000216 => x"E3500077",
000217 => x"1A00000C",
000218 => x"E3E03A0F",
000219 => x"E3A02050",
000220 => x"E5035F93",
000221 => x"E5032FAF",
000222 => x"E1A02003",
000223 => x"E5123FAF",
000224 => x"E3130002",
000225 => x"1AFFFFFC",
000226 => x"E5123FAF",
000227 => x"E2130080",
000228 => x"08BD8030",
000229 => x"E3E00002",
000230 => x"E8BD8030",
000231 => x"E3500072",
000232 => x"13E00003",
000233 => x"18BD8030",
000234 => x"E3813001",
000235 => x"E3E02A0F",
000236 => x"E3A01090",
000237 => x"E5023F93",
000238 => x"E5021FAF",
000239 => x"E5123FAF",
000240 => x"E3130002",
000241 => x"1AFFFFFC",
000242 => x"E5123FAF",
000243 => x"E3130080",
000244 => x"1AFFFFEF",
000245 => x"E3A03068",
000246 => x"E5023FAF",
000247 => x"E3E00A0F",
000248 => x"E5103FAF",
000249 => x"E3130002",
000250 => x"1AFFFFFC",
000251 => x"E5100F93",
000252 => x"E8BD8030",
000253 => x"E20000FF",
000254 => x"E350000F",
000255 => x"979FF100",
000256 => x"EA00000F",
000257 => x"000104C4",
000258 => x"000104BC",
000259 => x"000104B4",
000260 => x"000104AC",
000261 => x"000104A4",
000262 => x"0001049C",
000263 => x"00010494",
000264 => x"0001048C",
000265 => x"00010484",
000266 => x"0001047C",
000267 => x"00010474",
000268 => x"0001046C",
000269 => x"00010464",
000270 => x"0001045C",
000271 => x"00010454",
000272 => x"0001044C",
000273 => x"E3A00000",
000274 => x"E1A0F00E",
000275 => x"EE1F0F1F",
000276 => x"E1A0F00E",
000277 => x"EE1E0F1E",
000278 => x"E1A0F00E",
000279 => x"EE1D0F1D",
000280 => x"E1A0F00E",
000281 => x"EE1C0F1C",
000282 => x"E1A0F00E",
000283 => x"EE1B0F1B",
000284 => x"E1A0F00E",
000285 => x"EE1A0F1A",
000286 => x"E1A0F00E",
000287 => x"EE190F19",
000288 => x"E1A0F00E",
000289 => x"EE180F18",
000290 => x"E1A0F00E",
000291 => x"EE170F17",
000292 => x"E1A0F00E",
000293 => x"EE160F16",
000294 => x"E1A0F00E",
000295 => x"EE150F15",
000296 => x"E1A0F00E",
000297 => x"EE140F14",
000298 => x"E1A0F00E",
000299 => x"EE130F13",
000300 => x"E1A0F00E",
000301 => x"EE120F12",
000302 => x"E1A0F00E",
000303 => x"EE110F11",
000304 => x"E1A0F00E",
000305 => x"EE100F10",
000306 => x"E1A0F00E",
000307 => x"E20110FF",
000308 => x"E2411006",
000309 => x"E3510007",
000310 => x"979FF101",
000311 => x"EA000008",
000312 => x"00010508",
000313 => x"00010504",
000314 => x"00010504",
000315 => x"00010504",
000316 => x"00010504",
000317 => x"00010510",
000318 => x"00010518",
000319 => x"00010500",
000320 => x"EE0D0F1D",
000321 => x"E1A0F00E",
000322 => x"EE060F16",
000323 => x"E1A0F00E",
000324 => x"EE0B0F1B",
000325 => x"E1A0F00E",
000326 => x"EE0C0F1C",
000327 => x"E1A0F00E",
000328 => x"E92D4010",
000329 => x"E1A04000",
000330 => x"E5D00000",
000331 => x"E3500000",
000332 => x"1A000003",
000333 => x"EA000005",
000334 => x"E5F40001",
000335 => x"E3500000",
000336 => x"0A000002",
000337 => x"EBFFFF22",
000338 => x"E3500000",
000339 => x"CAFFFFF9",
000340 => x"E1A00004",
000341 => x"E8BD8010",
000342 => x"E92D4070",
000343 => x"E2514000",
000344 => x"E1A05000",
000345 => x"E20260FF",
000346 => x"D8BD8070",
000347 => x"EBFFFF12",
000348 => x"E3700001",
000349 => x"E20030FF",
000350 => x"0A000005",
000351 => x"E3560001",
000352 => x"E5C53000",
000353 => x"E1A00003",
000354 => x"E2855001",
000355 => x"0A000003",
000356 => x"E2444001",
000357 => x"E3540000",
000358 => x"CAFFFFF3",
000359 => x"E8BD8070",
000360 => x"EBFFFF0B",
000361 => x"EAFFFFF9",
000362 => x"E92D4030",
000363 => x"E2514000",
000364 => x"E1A05000",
000365 => x"D8BD8030",
000366 => x"E4D50001",
000367 => x"EBFFFF04",
000368 => x"E2544001",
000369 => x"1AFFFFFB",
000370 => x"E8BD8030",
000371 => x"E92D4010",
000372 => x"E20240FF",
000373 => x"E3540008",
000374 => x"83A04008",
000375 => x"8A000001",
000376 => x"E3540000",
000377 => x"03A04001",
000378 => x"E1A02001",
000379 => x"E1A0E004",
000380 => x"E1A0310E",
000381 => x"E35E0001",
000382 => x"E2433004",
000383 => x"E1A0C000",
000384 => x"81A0C330",
000385 => x"E24E3001",
000386 => x"E20CC00F",
000387 => x"E203E0FF",
000388 => x"E35C0009",
000389 => x"E28C3030",
000390 => x"828C3037",
000391 => x"E35E0000",
000392 => x"E4C23001",
000393 => x"1AFFFFF1",
000394 => x"E2443001",
000395 => x"E20330FF",
000396 => x"E0813003",
000397 => x"E5C3E001",
000398 => x"E8BD8010",
000399 => x"E92D4010",
000400 => x"E1A04000",
000401 => x"E3540007",
000402 => x"E3A01010",
000403 => x"E3A00001",
000404 => x"9A000001",
000405 => x"E3A00000",
000406 => x"E8BD8010",
000407 => x"EBFFFEE3",
000408 => x"E3A00006",
000409 => x"EBFFFEFB",
000410 => x"E3A00000",
000411 => x"EBFFFEEB",
000412 => x"E1A00584",
000413 => x"E8BD4010",
000414 => x"EAFFFEE8",
000415 => x"E0603280",
000416 => x"E0800103",
000417 => x"E0800100",
000418 => x"E1A00200",
000419 => x"E3500000",
000420 => x"D1A0F00E",
000421 => x"E1A00000",
000422 => x"E2500001",
000423 => x"1AFFFFFC",
000424 => x"E1A0F00E",
000425 => x"E212C0FF",
000426 => x"0A00000B",
000427 => x"E5D02000",
000428 => x"E5D13000",
000429 => x"E1520003",
000430 => x"0A000004",
000431 => x"EA000008",
000432 => x"E5F02001",
000433 => x"E5F13001",
000434 => x"E1520003",
000435 => x"1A000004",
000436 => x"E24C3001",
000437 => x"E213C0FF",
000438 => x"1AFFFFF8",
000439 => x"E3A00001",
000440 => x"E1A0F00E",
000441 => x"E3A00000",
000442 => x"E1A0F00E",
000443 => x"E92D4030",
000444 => x"E1A04081",
000445 => x"E3540000",
000446 => x"E1A05000",
000447 => x"D3A00000",
000448 => x"D8BD8030",
000449 => x"E3A00000",
000450 => x"E1A01000",
000451 => x"E7D12005",
000452 => x"E2423030",
000453 => x"E082C200",
000454 => x"E3530009",
000455 => x"E242E041",
000456 => x"924C0030",
000457 => x"9A000007",
000458 => x"E0823200",
000459 => x"E35E0005",
000460 => x"E242C061",
000461 => x"92430037",
000462 => x"9A000002",
000463 => x"E0823200",
000464 => x"E35C0005",
000465 => x"92430057",
000466 => x"E2811001",
000467 => x"E1510004",
000468 => x"1AFFFFED",
000469 => x"E8BD8030",
000470 => x"E5D03003",
000471 => x"E5D02002",
000472 => x"E5D01000",
000473 => x"E1833402",
000474 => x"E5D00001",
000475 => x"E1833C01",
000476 => x"E1830800",
000477 => x"E1A0F00E",
000478 => x"E92D45F0",
000479 => x"E3A00000",
000480 => x"E24DD00C",
000481 => x"EBFFFE56",
000482 => x"E3A0100D",
000483 => x"E3A000C3",
000484 => x"EBFFFF4D",
000485 => x"E3A00063",
000486 => x"EBFFFEBE",
000487 => x"E3A00006",
000488 => x"EBFFFF13",
000489 => x"E3A01006",
000490 => x"E3800008",
000491 => x"EBFFFF46",
000492 => x"E3A0000D",
000493 => x"EBFFFF0E",
000494 => x"E1A008A0",
000495 => x"E1E00000",
000496 => x"E200000F",
000497 => x"E3500001",
000498 => x"03A04030",
000499 => x"028DA007",
000500 => x"0A00001A",
000501 => x"E3500002",
000502 => x"0A000070",
000503 => x"E59F07EC",
000504 => x"EBFFFF4E",
000505 => x"E59F07E8",
000506 => x"EBFFFF4C",
000507 => x"E59F07E4",
000508 => x"EBFFFF4A",
000509 => x"E59F07E0",
000510 => x"EBFFFF48",
000511 => x"E59F07DC",
000512 => x"EBFFFF46",
000513 => x"E59F07D8",
000514 => x"EBFFFF44",
000515 => x"E59F07D4",
000516 => x"EBFFFF42",
000517 => x"E59F07D0",
000518 => x"EBFFFF40",
000519 => x"E59F07CC",
000520 => x"EBFFFF3E",
000521 => x"E59F07C8",
000522 => x"EBFFFF3C",
000523 => x"E59F07C4",
000524 => x"EBFFFF3A",
000525 => x"E28DA007",
000526 => x"EBFFFE5F",
000527 => x"E1A04000",
000528 => x"E3A0000D",
000529 => x"EBFFFEEA",
000530 => x"E3100801",
000531 => x"03A06001",
000532 => x"03A050A0",
000533 => x"1A000035",
000534 => x"E3A04000",
000535 => x"E59F0798",
000536 => x"EBFFFF2E",
000537 => x"E1A01005",
000538 => x"E1A02004",
000539 => x"E3A03002",
000540 => x"E3A00072",
000541 => x"E58D4000",
000542 => x"EBFFFE91",
000543 => x"E1A01005",
000544 => x"E5CD0007",
000545 => x"E3A02001",
000546 => x"E3A03002",
000547 => x"E3A00072",
000548 => x"E58D4000",
000549 => x"EBFFFE8A",
000550 => x"E3A02002",
000551 => x"E1A03002",
000552 => x"E5CD0008",
000553 => x"E1A01005",
000554 => x"E3A00072",
000555 => x"E58D4000",
000556 => x"EBFFFE83",
000557 => x"E3A03002",
000558 => x"E5CD0009",
000559 => x"E1A01005",
000560 => x"E3A00072",
000561 => x"E3A02003",
000562 => x"E58D4000",
000563 => x"EBFFFE7C",
000564 => x"E5DD3007",
000565 => x"E20000FF",
000566 => x"E3530053",
000567 => x"E5CD000A",
000568 => x"1A000002",
000569 => x"E5DD3008",
000570 => x"E353004D",
000571 => x"0A000062",
000572 => x"E59F0708",
000573 => x"EBFFFF09",
000574 => x"E3560000",
000575 => x"0AFFFFCD",
000576 => x"E59F06FC",
000577 => x"EBFFFF05",
000578 => x"E3A0100D",
000579 => x"E3A00000",
000580 => x"EBFFFEED",
000581 => x"E3A00006",
000582 => x"EBFFFEB5",
000583 => x"E3A01006",
000584 => x"E3C00008",
000585 => x"EBFFFEE8",
000586 => x"E3A0F000",
000587 => x"EAFFFFFE",
000588 => x"E3540034",
000589 => x"0A000028",
000590 => x"CA00001B",
000591 => x"E3540031",
000592 => x"0A000035",
000593 => x"DA000097",
000594 => x"E3540032",
000595 => x"0A0000A1",
000596 => x"E3540033",
000597 => x"1A000097",
000598 => x"E1A00004",
000599 => x"EBFFFE1C",
000600 => x"E59F06A0",
000601 => x"EBFFFEED",
000602 => x"E1A0000A",
000603 => x"E3A01002",
000604 => x"E3A02001",
000605 => x"EBFFFEF7",
000606 => x"E3A01002",
000607 => x"E1A0000A",
000608 => x"EBFFFF59",
000609 => x"E21010FF",
000610 => x"11A05001",
000611 => x"13A06000",
000612 => x"1AFFFFB0",
000613 => x"E59F0670",
000614 => x"EBFFFEE0",
000615 => x"EAFFFFA5",
000616 => x"E3A04033",
000617 => x"E28DA007",
000618 => x"EAFFFFA4",
000619 => x"E3540066",
000620 => x"0A00002A",
000621 => x"DA0000A5",
000622 => x"E3540068",
000623 => x"0A000107",
000624 => x"E3540072",
000625 => x"1A00007B",
000626 => x"E1A00004",
000627 => x"EBFFFE00",
000628 => x"E3A006FF",
000629 => x"E280F20F",
000630 => x"EAFFFFFE",
000631 => x"E1A00004",
000632 => x"EBFFFDFB",
000633 => x"E59F061C",
000634 => x"EBFFFECC",
000635 => x"E1A0000A",
000636 => x"E3A01002",
000637 => x"E3A02001",
000638 => x"EBFFFED6",
000639 => x"E1A0000A",
000640 => x"E3A01002",
000641 => x"EBFFFF38",
000642 => x"E21080FF",
000643 => x"1A00009C",
000644 => x"E59F05F8",
000645 => x"EBFFFEC1",
000646 => x"EAFFFF86",
000647 => x"E1A00004",
000648 => x"EBFFFDEB",
000649 => x"E59F05E8",
000650 => x"EBFFFEBC",
000651 => x"E1A0000A",
000652 => x"E3A01004",
000653 => x"E3A02000",
000654 => x"EBFFFEC6",
000655 => x"E5DD3007",
000656 => x"E3530053",
000657 => x"1A000002",
000658 => x"E5DD3008",
000659 => x"E353004D",
000660 => x"0A00010D",
000661 => x"E59F05BC",
000662 => x"EBFFFEB0",
000663 => x"EAFFFF75",
000664 => x"E1A00004",
000665 => x"EBFFFDDA",
000666 => x"E59F05AC",
000667 => x"EBFFFEAB",
000668 => x"E59F05A8",
000669 => x"EBFFFEA9",
000670 => x"EAFFFF6E",
000671 => x"E5DD3009",
000672 => x"E3530042",
000673 => x"1AFFFF99",
000674 => x"E3500052",
000675 => x"1AFFFF97",
000676 => x"E1A01005",
000677 => x"E3A02004",
000678 => x"E2433040",
000679 => x"E2800020",
000680 => x"E58D4000",
000681 => x"EBFFFE06",
000682 => x"E1A01005",
000683 => x"E5CD0007",
000684 => x"E3A02005",
000685 => x"E3A03002",
000686 => x"E3A00072",
000687 => x"E58D4000",
000688 => x"EBFFFDFF",
000689 => x"E1A01005",
000690 => x"E5CD0008",
000691 => x"E3A02006",
000692 => x"E3A03002",
000693 => x"E3A00072",
000694 => x"E58D4000",
000695 => x"EBFFFDF8",
000696 => x"E1A01005",
000697 => x"E5CD0009",
000698 => x"E3A02007",
000699 => x"E3A03002",
000700 => x"E3A00072",
000701 => x"E58D4000",
000702 => x"EBFFFDF1",
000703 => x"E5CD000A",
000704 => x"E1A0000A",
000705 => x"EBFFFF13",
000706 => x"E2907004",
000707 => x"0A000022",
000708 => x"E1A06004",
000709 => x"E2842008",
000710 => x"E1A01005",
000711 => x"E3A03002",
000712 => x"E3A00072",
000713 => x"E58D6000",
000714 => x"EBFFFDE5",
000715 => x"E2842009",
000716 => x"E5CD0007",
000717 => x"E1A01005",
000718 => x"E3A03002",
000719 => x"E3A00072",
000720 => x"E58D6000",
000721 => x"EBFFFDDE",
000722 => x"E284200A",
000723 => x"E5CD0008",
000724 => x"E1A01005",
000725 => x"E3A03002",
000726 => x"E3A00072",
000727 => x"E58D6000",
000728 => x"EBFFFDD7",
000729 => x"E284200B",
000730 => x"E5CD0009",
000731 => x"E1A01005",
000732 => x"E3A03002",
000733 => x"E3A00072",
000734 => x"E58D6000",
000735 => x"EBFFFDD0",
000736 => x"E5CD000A",
000737 => x"E1A0000A",
000738 => x"EBFFFEF2",
000739 => x"E4840004",
000740 => x"E1540007",
000741 => x"13540902",
000742 => x"3AFFFFDD",
000743 => x"E59F0480",
000744 => x"EBFFFE5E",
000745 => x"EAFFFF55",
000746 => x"E3740001",
000747 => x"0AFFFF21",
000748 => x"E3540030",
000749 => x"0A000004",
000750 => x"E20400FF",
000751 => x"EBFFFD84",
000752 => x"E59F0460",
000753 => x"EBFFFE55",
000754 => x"EAFFFF1A",
000755 => x"E1A00004",
000756 => x"EBFFFD7F",
000757 => x"EAFFFF49",
000758 => x"E1A00004",
000759 => x"EBFFFD7C",
000760 => x"E59F0444",
000761 => x"EBFFFE4D",
000762 => x"EBFFFD73",
000763 => x"E3700001",
000764 => x"0AFFFFFC",
000765 => x"EBFFFD70",
000766 => x"E3700001",
000767 => x"1AFFFFFC",
000768 => x"E3A05000",
000769 => x"EA000001",
000770 => x"E3550902",
000771 => x"0A00000C",
000772 => x"E5954000",
000773 => x"E1A00C24",
000774 => x"EBFFFD6D",
000775 => x"E1A00824",
000776 => x"EBFFFD6B",
000777 => x"E1A00424",
000778 => x"EBFFFD69",
000779 => x"E1A00004",
000780 => x"EBFFFD67",
000781 => x"EBFFFD60",
000782 => x"E3700001",
000783 => x"E2855004",
000784 => x"0AFFFFF0",
000785 => x"E59F03E4",
000786 => x"EBFFFE34",
000787 => x"EAFFFEF9",
000788 => x"E3540035",
000789 => x"0A0000A9",
000790 => x"E3540061",
000791 => x"1AFFFFD5",
000792 => x"E1A00004",
000793 => x"EBFFFD5A",
000794 => x"E59F03C4",
000795 => x"EBFFFE2B",
000796 => x"E59F03C0",
000797 => x"EBFFFE29",
000798 => x"E59F03BC",
000799 => x"EBFFFE27",
000800 => x"EAFFFEEC",
000801 => x"E59F03B4",
000802 => x"EBFFFE24",
000803 => x"E1A0000A",
000804 => x"E3A01004",
000805 => x"E3A02000",
000806 => x"EBFFFE2E",
000807 => x"E5DD3007",
000808 => x"E3530053",
000809 => x"1A000002",
000810 => x"E5DD2008",
000811 => x"E352004D",
000812 => x"0A000004",
000813 => x"E59F0388",
000814 => x"EBFFFE18",
000815 => x"E59F0384",
000816 => x"EBFFFE16",
000817 => x"EAFFFEDB",
000818 => x"E5DD1009",
000819 => x"E3510042",
000820 => x"1AFFFFF7",
000821 => x"E5DD000A",
000822 => x"E3500052",
000823 => x"1AFFFFF4",
000824 => x"E3A04000",
000825 => x"E5C43000",
000826 => x"E1A00000",
000827 => x"E5C42001",
000828 => x"E1A00000",
000829 => x"E5C41002",
000830 => x"E1A00000",
000831 => x"E5C40003",
000832 => x"E1A00000",
000833 => x"E241103E",
000834 => x"E1A0000A",
000835 => x"E1A02004",
000836 => x"EBFFFE10",
000837 => x"E5DD3007",
000838 => x"E5C43004",
000839 => x"E5DD2008",
000840 => x"E5C42005",
000841 => x"E5DD3009",
000842 => x"E5C43006",
000843 => x"E5DD200A",
000844 => x"E1A0000A",
000845 => x"E5C42007",
000846 => x"EBFFFE86",
000847 => x"E3A03CFF",
000848 => x"E28330FC",
000849 => x"E1500003",
000850 => x"E1A05000",
000851 => x"8A000095",
000852 => x"E3700004",
000853 => x"12844008",
000854 => x"1280600B",
000855 => x"0A000006",
000856 => x"EBFFFD15",
000857 => x"E3700001",
000858 => x"0AFFFFFC",
000859 => x"E1560004",
000860 => x"E5C40000",
000861 => x"E2844001",
000862 => x"1AFFFFF8",
000863 => x"E59F02C8",
000864 => x"EBFFFDE6",
000865 => x"E59F02C4",
000866 => x"EBFFFDE4",
000867 => x"E375000C",
000868 => x"0A00000F",
000869 => x"E3A04000",
000870 => x"E285700C",
000871 => x"E1A06004",
000872 => x"E5D45000",
000873 => x"E3A00077",
000874 => x"E1A01008",
000875 => x"E1A02006",
000876 => x"E3A03002",
000877 => x"E58D5000",
000878 => x"EBFFFD41",
000879 => x"E3500000",
000880 => x"1AFFFFF7",
000881 => x"E2844001",
000882 => x"E1540007",
000883 => x"E1A06004",
000884 => x"1AFFFFF2",
000885 => x"E59F0278",
000886 => x"EBFFFDD0",
000887 => x"EAFFFFB6",
000888 => x"E1A00004",
000889 => x"EBFFFCFA",
000890 => x"E59F0268",
000891 => x"EBFFFDCB",
000892 => x"E59F0264",
000893 => x"EBFFFDC9",
000894 => x"E59F0260",
000895 => x"EBFFFDC7",
000896 => x"E59F025C",
000897 => x"EBFFFDC5",
000898 => x"E59F0258",
000899 => x"EBFFFDC3",
000900 => x"E59F0254",
000901 => x"EBFFFDC1",
000902 => x"E59F0250",
000903 => x"EBFFFDBF",
000904 => x"E59F024C",
000905 => x"EBFFFDBD",
000906 => x"E59F0248",
000907 => x"EBFFFDBB",
000908 => x"E59F0244",
000909 => x"EBFFFDB9",
000910 => x"E59F0240",
000911 => x"EBFFFDB7",
000912 => x"E59F023C",
000913 => x"EBFFFDB5",
000914 => x"E59F0238",
000915 => x"EBFFFDB3",
000916 => x"E59F0234",
000917 => x"EBFFFDB1",
000918 => x"E59F0230",
000919 => x"EBFFFDAF",
000920 => x"E59F022C",
000921 => x"EBFFFDAD",
000922 => x"E59F0228",
000923 => x"EBFFFDAB",
000924 => x"E59F0224",
000925 => x"EBFFFDA9",
000926 => x"E59F0220",
000927 => x"EBFFFDA7",
000928 => x"E59F021C",
000929 => x"EBFFFDA5",
000930 => x"EAFFFE6A",
000931 => x"E5DD3009",
000932 => x"E3530042",
000933 => x"1AFFFEEE",
000934 => x"E5DD300A",
000935 => x"E3530052",
000936 => x"1AFFFEEB",
000937 => x"E3A01004",
000938 => x"E3A02000",
000939 => x"E1A0000A",
000940 => x"EBFFFDA8",
000941 => x"E1A0000A",
000942 => x"EBFFFE26",
000943 => x"E3A03C7F",
000944 => x"E28330F8",
000945 => x"E1500003",
000946 => x"8A000036",
000947 => x"E2905004",
000948 => x"0AFFFE8A",
000949 => x"E3A04000",
000950 => x"E3A01004",
000951 => x"E3A02000",
000952 => x"E1A0000A",
000953 => x"EBFFFD9B",
000954 => x"E1A0000A",
000955 => x"EBFFFE19",
000956 => x"E4840004",
000957 => x"E1550004",
000958 => x"1AFFFFF6",
000959 => x"EAFFFE7F",
000960 => x"E1A00004",
000961 => x"EBFFFCB2",
000962 => x"E59F0198",
000963 => x"EBFFFD83",
000964 => x"E1A0000A",
000965 => x"E3A01002",
000966 => x"E3A02001",
000967 => x"EBFFFD8D",
000968 => x"E1A0000A",
000969 => x"E3A01002",
000970 => x"EBFFFDEF",
000971 => x"E21060FF",
000972 => x"0AFFFE97",
000973 => x"E59F0170",
000974 => x"EBFFFD78",
000975 => x"E59F016C",
000976 => x"EBFFFD76",
000977 => x"EBFFFC9C",
000978 => x"E3700001",
000979 => x"0AFFFFFC",
000980 => x"EBFFFC99",
000981 => x"E3700001",
000982 => x"1AFFFFFC",
000983 => x"E3A05000",
000984 => x"EA000001",
000985 => x"E3540000",
000986 => x"AA000011",
000987 => x"E3A0C000",
000988 => x"E1A02005",
000989 => x"E1A01006",
000990 => x"E3A03002",
000991 => x"E3A00072",
000992 => x"E58DC000",
000993 => x"EBFFFCCE",
000994 => x"E1A04000",
000995 => x"EBFFFC8A",
000996 => x"E3700001",
000997 => x"E1A00004",
000998 => x"0AFFFFF1",
000999 => x"E59F0110",
001000 => x"EBFFFD5E",
001001 => x"EAFFFF26",
001002 => x"E59F0108",
001003 => x"EBFFFD5B",
001004 => x"EAFFFE20",
001005 => x"EBFFFC86",
001006 => x"E3A03801",
001007 => x"E2855001",
001008 => x"E2433001",
001009 => x"E1550003",
001010 => x"1AFFFFE7",
001011 => x"EAFFFF1C",
001012 => x"000110DC",
001013 => x"00011128",
001014 => x"00011170",
001015 => x"000111B8",
001016 => x"00011200",
001017 => x"00011248",
001018 => x"00011290",
001019 => x"000112FC",
001020 => x"00011334",
001021 => x"00011398",
001022 => x"000113FC",
001023 => x"000115D4",
001024 => x"00011638",
001025 => x"00011D3C",
001026 => x"00011578",
001027 => x"000115B4",
001028 => x"00011664",
001029 => x"0001144C",
001030 => x"000114E4",
001031 => x"00011CC0",
001032 => x"00011CF0",
001033 => x"00011624",
001034 => x"00011D18",
001035 => x"0001150C",
001036 => x"00011554",
001037 => x"00011814",
001038 => x"00011848",
001039 => x"000118B4",
001040 => x"00011684",
001041 => x"0001172C",
001042 => x"00011D0C",
001043 => x"000116E4",
001044 => x"000116FC",
001045 => x"0001171C",
001046 => x"000118F8",
001047 => x"00011914",
001048 => x"00011934",
001049 => x"00011974",
001050 => x"000119A8",
001051 => x"000119E4",
001052 => x"00011A20",
001053 => x"00011A44",
001054 => x"00011A80",
001055 => x"00011A9C",
001056 => x"00011AB4",
001057 => x"00011AFC",
001058 => x"00011B3C",
001059 => x"00011B74",
001060 => x"00011B98",
001061 => x"00011BDC",
001062 => x"00011C1C",
001063 => x"00011C48",
001064 => x"00011C74",
001065 => x"00011C98",
001066 => x"00011750",
001067 => x"0001178C",
001068 => x"000117CC",
001069 => x"00011D60",
001070 => x"000114C0",
001071 => x"E10F3000",
001072 => x"E3C330C0",
001073 => x"E129F003",
001074 => x"E1A0F00E",
001075 => x"E10F3000",
001076 => x"E38330C0",
001077 => x"E129F003",
001078 => x"E1A0F00E",
001079 => x"0D0A0D0A",
001080 => x"0D0A2B2D",
001081 => x"2D2D2D2D",
001082 => x"2D2D2D2D",
001083 => x"2D2D2D2D",
001084 => x"2D2D2D2D",
001085 => x"2D2D2D2D",
001086 => x"2D2D2D2D",
001087 => x"2D2D2D2D",
001088 => x"2D2D2D2D",
001089 => x"2D2D2D2D",
001090 => x"2D2D2D2D",
001091 => x"2D2D2D2D",
001092 => x"2D2D2D2D",
001093 => x"2D2D2D2D",
001094 => x"2D2D2D2D",
001095 => x"2D2D2D2D",
001096 => x"2D2D2D2B",
001097 => x"0D0A0000",
001098 => x"7C202020",
001099 => x"203C3C3C",
001100 => x"2053544F",
001101 => x"524D2043",
001102 => x"6F726520",
001103 => x"50726F63",
001104 => x"6573736F",
001105 => x"72205379",
001106 => x"7374656D",
001107 => x"202D2042",
001108 => x"79205374",
001109 => x"65706861",
001110 => x"6E204E6F",
001111 => x"6C74696E",
001112 => x"67203E3E",
001113 => x"3E202020",
001114 => x"207C0D0A",
001115 => x"00000000",
001116 => x"2B2D2D2D",
001117 => x"2D2D2D2D",
001118 => x"2D2D2D2D",
001119 => x"2D2D2D2D",
001120 => x"2D2D2D2D",
001121 => x"2D2D2D2D",
001122 => x"2D2D2D2D",
001123 => x"2D2D2D2D",
001124 => x"2D2D2D2D",
001125 => x"2D2D2D2D",
001126 => x"2D2D2D2D",
001127 => x"2D2D2D2D",
001128 => x"2D2D2D2D",
001129 => x"2D2D2D2D",
001130 => x"2D2D2D2D",
001131 => x"2D2D2D2D",
001132 => x"2D2B0D0A",
001133 => x"00000000",
001134 => x"7C202020",
001135 => x"20202020",
001136 => x"2020426F",
001137 => x"6F746C6F",
001138 => x"61646572",
001139 => x"20666F72",
001140 => x"2053544F",
001141 => x"524D2053",
001142 => x"6F432020",
001143 => x"20566572",
001144 => x"73696F6E",
001145 => x"3A203230",
001146 => x"31323035",
001147 => x"32342D44",
001148 => x"20202020",
001149 => x"20202020",
001150 => x"207C0D0A",
001151 => x"00000000",
001152 => x"7C202020",
001153 => x"20202020",
001154 => x"20202020",
001155 => x"20202020",
001156 => x"436F6E74",
001157 => x"6163743A",
001158 => x"2073746E",
001159 => x"6F6C7469",
001160 => x"6E674067",
001161 => x"6F6F676C",
001162 => x"656D6169",
001163 => x"6C2E636F",
001164 => x"6D202020",
001165 => x"20202020",
001166 => x"20202020",
001167 => x"20202020",
001168 => x"207C0D0A",
001169 => x"00000000",
001170 => x"2B2D2D2D",
001171 => x"2D2D2D2D",
001172 => x"2D2D2D2D",
001173 => x"2D2D2D2D",
001174 => x"2D2D2D2D",
001175 => x"2D2D2D2D",
001176 => x"2D2D2D2D",
001177 => x"2D2D2D2D",
001178 => x"2D2D2D2D",
001179 => x"2D2D2D2D",
001180 => x"2D2D2D2D",
001181 => x"2D2D2D2D",
001182 => x"2D2D2D2D",
001183 => x"2D2D2D2D",
001184 => x"2D2D2D2D",
001185 => x"2D2D2D2D",
001186 => x"2D2B0D0A",
001187 => x"0D0A0000",
001188 => x"203C2057",
001189 => x"656C636F",
001190 => x"6D652074",
001191 => x"6F207468",
001192 => x"65205354",
001193 => x"4F524D20",
001194 => x"536F4320",
001195 => x"626F6F74",
001196 => x"6C6F6164",
001197 => x"65722063",
001198 => x"6F6E736F",
001199 => x"6C652120",
001200 => x"3E0D0A20",
001201 => x"3C205365",
001202 => x"6C656374",
001203 => x"20616E20",
001204 => x"6F706572",
001205 => x"6174696F",
001206 => x"6E206672",
001207 => x"6F6D2074",
001208 => x"6865206D",
001209 => x"656E7520",
001210 => x"62656C6F",
001211 => x"77206F72",
001212 => x"20707265",
001213 => x"7373203E",
001214 => x"0D0A0000",
001215 => x"203C2074",
001216 => x"68652062",
001217 => x"6F6F7420",
001218 => x"6B657920",
001219 => x"666F7220",
001220 => x"696D6D65",
001221 => x"64696174",
001222 => x"65206170",
001223 => x"706C6963",
001224 => x"6174696F",
001225 => x"6E207374",
001226 => x"6172742E",
001227 => x"203E0D0A",
001228 => x"0D0A0000",
001229 => x"2030202D",
001230 => x"20626F6F",
001231 => x"74206672",
001232 => x"6F6D2063",
001233 => x"6F726520",
001234 => x"52414D20",
001235 => x"28737461",
001236 => x"72742061",
001237 => x"70706C69",
001238 => x"63617469",
001239 => x"6F6E290D",
001240 => x"0A203120",
001241 => x"2D207072",
001242 => x"6F677261",
001243 => x"6D20636F",
001244 => x"72652052",
001245 => x"414D2076",
001246 => x"69612055",
001247 => x"4152545F",
001248 => x"300D0A20",
001249 => x"32202D20",
001250 => x"636F7265",
001251 => x"2052414D",
001252 => x"2064756D",
001253 => x"700D0A00",
001254 => x"2033202D",
001255 => x"20626F6F",
001256 => x"74206672",
001257 => x"6F6D2049",
001258 => x"32432045",
001259 => x"4550524F",
001260 => x"4D0D0A20",
001261 => x"34202D20",
001262 => x"70726F67",
001263 => x"72616D20",
001264 => x"49324320",
001265 => x"45455052",
001266 => x"4F4D2076",
001267 => x"69612055",
001268 => x"4152545F",
001269 => x"300D0A20",
001270 => x"35202D20",
001271 => x"73686F77",
001272 => x"20636F6E",
001273 => x"74656E74",
001274 => x"206F6620",
001275 => x"49324320",
001276 => x"45455052",
001277 => x"4F4D0D0A",
001278 => x"00000000",
001279 => x"2061202D",
001280 => x"20617574",
001281 => x"6F6D6174",
001282 => x"69632062",
001283 => x"6F6F7420",
001284 => x"636F6E66",
001285 => x"69677572",
001286 => x"6174696F",
001287 => x"6E0D0A20",
001288 => x"68202D20",
001289 => x"68656C70",
001290 => x"0D0A2072",
001291 => x"202D2072",
001292 => x"65737461",
001293 => x"72742073",
001294 => x"79737465",
001295 => x"6D0D0A0D",
001296 => x"0A53656C",
001297 => x"6563743A",
001298 => x"20000000",
001299 => x"0D0A0D0A",
001300 => x"4170706C",
001301 => x"69636174",
001302 => x"696F6E20",
001303 => x"77696C6C",
001304 => x"20737461",
001305 => x"72742061",
001306 => x"75746F6D",
001307 => x"61746963",
001308 => x"616C6C79",
001309 => x"20616674",
001310 => x"65722064",
001311 => x"6F776E6C",
001312 => x"6F61642E",
001313 => x"0D0A2D3E",
001314 => x"20576169",
001315 => x"74696E67",
001316 => x"20666F72",
001317 => x"20277374",
001318 => x"6F726D5F",
001319 => x"70726F67",
001320 => x"72616D2E",
001321 => x"62696E27",
001322 => x"20696E20",
001323 => x"62797465",
001324 => x"2D737472",
001325 => x"65616D20",
001326 => x"6D6F6465",
001327 => x"2E2E2E00",
001328 => x"20455252",
001329 => x"4F522120",
001330 => x"50726F67",
001331 => x"72616D20",
001332 => x"66696C65",
001333 => x"20746F6F",
001334 => x"20626967",
001335 => x"210D0A0D",
001336 => x"0A000000",
001337 => x"20496E76",
001338 => x"616C6964",
001339 => x"2070726F",
001340 => x"6772616D",
001341 => x"6D696E67",
001342 => x"2066696C",
001343 => x"65210D0A",
001344 => x"0D0A5365",
001345 => x"6C656374",
001346 => x"3A200000",
001347 => x"0D0A0D0A",
001348 => x"41626F72",
001349 => x"74206475",
001350 => x"6D70696E",
001351 => x"67206279",
001352 => x"20707265",
001353 => x"7373696E",
001354 => x"6720616E",
001355 => x"79206B65",
001356 => x"792E0D0A",
001357 => x"50726573",
001358 => x"7320616E",
001359 => x"79206B65",
001360 => x"7920746F",
001361 => x"20636F6E",
001362 => x"74696E75",
001363 => x"652E0D0A",
001364 => x"0D0A0000",
001365 => x"0D0A0D0A",
001366 => x"44756D70",
001367 => x"696E6720",
001368 => x"636F6D70",
001369 => x"6C657465",
001370 => x"642E0D0A",
001371 => x"0D0A5365",
001372 => x"6C656374",
001373 => x"3A200000",
001374 => x"0D0A0D0A",
001375 => x"456E7465",
001376 => x"72206465",
001377 => x"76696365",
001378 => x"20616464",
001379 => x"72657373",
001380 => x"20283278",
001381 => x"20686578",
001382 => x"5F636861",
001383 => x"72732C20",
001384 => x"73657420",
001385 => x"4C534220",
001386 => x"746F2027",
001387 => x"3027293A",
001388 => x"20000000",
001389 => x"20496E76",
001390 => x"616C6964",
001391 => x"20616464",
001392 => x"72657373",
001393 => x"210D0A0D",
001394 => x"0A53656C",
001395 => x"6563743A",
001396 => x"20000000",
001397 => x"0D0A4170",
001398 => x"706C6963",
001399 => x"6174696F",
001400 => x"6E207769",
001401 => x"6C6C2073",
001402 => x"74617274",
001403 => x"20617574",
001404 => x"6F6D6174",
001405 => x"6963616C",
001406 => x"6C792061",
001407 => x"66746572",
001408 => x"2075706C",
001409 => x"6F61642E",
001410 => x"0D0A2D3E",
001411 => x"204C6F61",
001412 => x"64696E67",
001413 => x"20626F6F",
001414 => x"7420696D",
001415 => x"6167652E",
001416 => x"2E2E0000",
001417 => x"2055706C",
001418 => x"6F616420",
001419 => x"636F6D70",
001420 => x"6C657465",
001421 => x"0D0A0000",
001422 => x"20496E76",
001423 => x"616C6964",
001424 => x"20626F6F",
001425 => x"74206465",
001426 => x"76696365",
001427 => x"206F7220",
001428 => x"66696C65",
001429 => x"210D0A0D",
001430 => x"0A53656C",
001431 => x"6563743A",
001432 => x"20000000",
001433 => x"0D0A496E",
001434 => x"76616C69",
001435 => x"64206164",
001436 => x"64726573",
001437 => x"73210D0A",
001438 => x"0D0A5365",
001439 => x"6C656374",
001440 => x"3A200000",
001441 => x"0D0A4461",
001442 => x"74612077",
001443 => x"696C6C20",
001444 => x"6F766572",
001445 => x"77726974",
001446 => x"65205241",
001447 => x"4D20636F",
001448 => x"6E74656E",
001449 => x"74210D0A",
001450 => x"2D3E2057",
001451 => x"61697469",
001452 => x"6E672066",
001453 => x"6F722027",
001454 => x"73746F72",
001455 => x"6D5F7072",
001456 => x"6F677261",
001457 => x"6D2E6269",
001458 => x"6E272069",
001459 => x"6E206279",
001460 => x"74652D73",
001461 => x"74726561",
001462 => x"6D206D6F",
001463 => x"64652E2E",
001464 => x"2E000000",
001465 => x"20446F77",
001466 => x"6E6C6F61",
001467 => x"6420636F",
001468 => x"6D706C65",
001469 => x"7465640D",
001470 => x"0A000000",
001471 => x"57726974",
001472 => x"696E6720",
001473 => x"62756666",
001474 => x"65722074",
001475 => x"6F206932",
001476 => x"63204545",
001477 => x"50524F4D",
001478 => x"2E2E2E00",
001479 => x"20436F6D",
001480 => x"706C6574",
001481 => x"65640D0A",
001482 => x"0D0A0000",
001483 => x"20496E76",
001484 => x"616C6964",
001485 => x"20626F6F",
001486 => x"74206465",
001487 => x"76696365",
001488 => x"206F7220",
001489 => x"66696C65",
001490 => x"210D0A0D",
001491 => x"0A000000",
001492 => x"0D0A0D0A",
001493 => x"456E7465",
001494 => x"72206465",
001495 => x"76696365",
001496 => x"20616464",
001497 => x"72657373",
001498 => x"20283220",
001499 => x"6865782D",
001500 => x"63686172",
001501 => x"732C2073",
001502 => x"6574204C",
001503 => x"53422074",
001504 => x"6F202730",
001505 => x"27293A20",
001506 => x"00000000",
001507 => x"0D0A0D0A",
001508 => x"41626F72",
001509 => x"74206475",
001510 => x"6D70696E",
001511 => x"67206279",
001512 => x"20707265",
001513 => x"7373696E",
001514 => x"6720616E",
001515 => x"79206B65",
001516 => x"792E2049",
001517 => x"66206E6F",
001518 => x"20646174",
001519 => x"61206973",
001520 => x"2073686F",
001521 => x"776E2C0D",
001522 => x"0A000000",
001523 => x"74686520",
001524 => x"73656C65",
001525 => x"63746564",
001526 => x"20646576",
001527 => x"69636520",
001528 => x"6973206E",
001529 => x"6F742072",
001530 => x"6573706F",
001531 => x"6E64696E",
001532 => x"672E2050",
001533 => x"72657373",
001534 => x"20616E79",
001535 => x"206B6579",
001536 => x"20746F20",
001537 => x"636F6E74",
001538 => x"696E7565",
001539 => x"2E0D0A0D",
001540 => x"0A000000",
001541 => x"0D0A0D0A",
001542 => x"4175746F",
001543 => x"6D617469",
001544 => x"6320626F",
001545 => x"6F742063",
001546 => x"6F6E6669",
001547 => x"67757261",
001548 => x"74696F6E",
001549 => x"20666F72",
001550 => x"20706F77",
001551 => x"65722D75",
001552 => x"703A0D0A",
001553 => x"00000000",
001554 => x"5B333231",
001555 => x"305D2063",
001556 => x"6F6E6669",
001557 => x"67757261",
001558 => x"74696F6E",
001559 => x"20444950",
001560 => x"20737769",
001561 => x"7463680D",
001562 => x"0A203030",
001563 => x"3030202D",
001564 => x"20537461",
001565 => x"72742062",
001566 => x"6F6F746C",
001567 => x"6F616465",
001568 => x"7220636F",
001569 => x"6E736F6C",
001570 => x"650D0A20",
001571 => x"30303031",
001572 => x"202D2041",
001573 => x"75746F6D",
001574 => x"61746963",
001575 => x"20626F6F",
001576 => x"74206672",
001577 => x"6F6D2063",
001578 => x"6F726520",
001579 => x"52414D0D",
001580 => x"0A000000",
001581 => x"20303031",
001582 => x"30202D20",
001583 => x"4175746F",
001584 => x"6D617469",
001585 => x"6320626F",
001586 => x"6F742066",
001587 => x"726F6D20",
001588 => x"49324320",
001589 => x"45455052",
001590 => x"4F4D2028",
001591 => x"41646472",
001592 => x"65737320",
001593 => x"30784130",
001594 => x"290D0A0D",
001595 => x"0A53656C",
001596 => x"6563743A",
001597 => x"20000000",
001598 => x"0D0A0D0A",
001599 => x"53544F52",
001600 => x"4D20536F",
001601 => x"4320626F",
001602 => x"6F746C6F",
001603 => x"61646572",
001604 => x"0D0A0000",
001605 => x"2730273A",
001606 => x"20457865",
001607 => x"63757465",
001608 => x"2070726F",
001609 => x"6772616D",
001610 => x"20696E20",
001611 => x"52414D2E",
001612 => x"0D0A0000",
001613 => x"2731273A",
001614 => x"20577269",
001615 => x"74652027",
001616 => x"73746F72",
001617 => x"6D5F7072",
001618 => x"6F677261",
001619 => x"6D2E6269",
001620 => x"6E272074",
001621 => x"6F207468",
001622 => x"6520636F",
001623 => x"72652773",
001624 => x"2052414D",
001625 => x"20766961",
001626 => x"20554152",
001627 => x"542E0D0A",
001628 => x"00000000",
001629 => x"2732273A",
001630 => x"20507269",
001631 => x"6E742063",
001632 => x"75727265",
001633 => x"6E742063",
001634 => x"6F6E7465",
001635 => x"6E74206F",
001636 => x"6620636F",
001637 => x"6D706C65",
001638 => x"74652063",
001639 => x"6F726520",
001640 => x"52414D2E",
001641 => x"0D0A0000",
001642 => x"2733273A",
001643 => x"204C6F61",
001644 => x"6420626F",
001645 => x"6F742069",
001646 => x"6D616765",
001647 => x"2066726F",
001648 => x"6D204545",
001649 => x"50524F4D",
001650 => x"20616E64",
001651 => x"20737461",
001652 => x"72742061",
001653 => x"70706C69",
001654 => x"63617469",
001655 => x"6F6E2E0D",
001656 => x"0A000000",
001657 => x"2734273A",
001658 => x"20577269",
001659 => x"74652027",
001660 => x"73746F72",
001661 => x"6D5F7072",
001662 => x"6F677261",
001663 => x"6D2E6269",
001664 => x"6E272074",
001665 => x"6F204932",
001666 => x"43204545",
001667 => x"50524F4D",
001668 => x"20766961",
001669 => x"20554152",
001670 => x"542E0D0A",
001671 => x"00000000",
001672 => x"2735273A",
001673 => x"20507269",
001674 => x"6E742063",
001675 => x"6F6E7465",
001676 => x"6E74206F",
001677 => x"66204932",
001678 => x"43204545",
001679 => x"50524F4D",
001680 => x"2E0D0A00",
001681 => x"2761273A",
001682 => x"2053686F",
001683 => x"77204449",
001684 => x"50207377",
001685 => x"69746368",
001686 => x"20636F6E",
001687 => x"66696775",
001688 => x"72617469",
001689 => x"6F6E7320",
001690 => x"666F7220",
001691 => x"6175746F",
001692 => x"6D617469",
001693 => x"6320626F",
001694 => x"6F742E0D",
001695 => x"0A000000",
001696 => x"2768273A",
001697 => x"2053686F",
001698 => x"77207468",
001699 => x"69732073",
001700 => x"63726565",
001701 => x"6E2E0D0A",
001702 => x"00000000",
001703 => x"2772273A",
001704 => x"20526573",
001705 => x"65742073",
001706 => x"79737465",
001707 => x"6D2E0D0A",
001708 => x"0D0A0000",
001709 => x"426F6F74",
001710 => x"20454550",
001711 => x"524F4D3A",
001712 => x"20323478",
001713 => x"786E6E6E",
001714 => x"20286C69",
001715 => x"6B652032",
001716 => x"34414136",
001717 => x"34292C20",
001718 => x"37206269",
001719 => x"74206164",
001720 => x"64726573",
001721 => x"73202B20",
001722 => x"646F6E74",
001723 => x"2D636172",
001724 => x"65206269",
001725 => x"742C0D0A",
001726 => x"00000000",
001727 => x"636F6E6E",
001728 => x"65637465",
001729 => x"6420746F",
001730 => x"20493243",
001731 => x"5F434F4E",
001732 => x"54524F4C",
001733 => x"4C45525F",
001734 => x"302C206F",
001735 => x"70657261",
001736 => x"74696E67",
001737 => x"20667265",
001738 => x"7175656E",
001739 => x"63792069",
001740 => x"73203130",
001741 => x"306B487A",
001742 => x"2C0D0A00",
001743 => x"6D617869",
001744 => x"6D756D20",
001745 => x"45455052",
001746 => x"4F4D2073",
001747 => x"697A6520",
001748 => x"3D203635",
001749 => x"35333620",
001750 => x"62797465",
001751 => x"203D3E20",
001752 => x"31362062",
001753 => x"69742061",
001754 => x"64647265",
001755 => x"73736573",
001756 => x"2C0D0A00",
001757 => x"66697865",
001758 => x"6420626F",
001759 => x"6F742064",
001760 => x"65766963",
001761 => x"65206164",
001762 => x"64726573",
001763 => x"733A2030",
001764 => x"7841300D",
001765 => x"0A0D0A00",
001766 => x"5465726D",
001767 => x"696E616C",
001768 => x"20736574",
001769 => x"75703A20",
001770 => x"39363030",
001771 => x"20626175",
001772 => x"642C2038",
001773 => x"20646174",
001774 => x"61206269",
001775 => x"74732C20",
001776 => x"6E6F2070",
001777 => x"61726974",
001778 => x"792C2031",
001779 => x"2073746F",
001780 => x"70206269",
001781 => x"740D0A0D",
001782 => x"0A000000",
001783 => x"466F7220",
001784 => x"6D6F7265",
001785 => x"20696E66",
001786 => x"6F726D61",
001787 => x"74696F6E",
001788 => x"20736565",
001789 => x"20746865",
001790 => x"2053544F",
001791 => x"524D2043",
001792 => x"6F726520",
001793 => x"2F205354",
001794 => x"4F524D20",
001795 => x"536F4320",
001796 => x"64617461",
001797 => x"73686565",
001798 => x"740D0A00",
001799 => x"68747470",
001800 => x"3A2F2F6F",
001801 => x"70656E63",
001802 => x"6F726573",
001803 => x"2E6F7267",
001804 => x"2F70726F",
001805 => x"6A656374",
001806 => x"2C73746F",
001807 => x"726D5F63",
001808 => x"6F72650D",
001809 => x"0A000000",
001810 => x"68747470",
001811 => x"3A2F2F6F",
001812 => x"70656E63",
001813 => x"6F726573",
001814 => x"2E6F7267",
001815 => x"2F70726F",
001816 => x"6A656374",
001817 => x"2C73746F",
001818 => x"726D5F73",
001819 => x"6F630D0A",
001820 => x"00000000",
001821 => x"436F6E74",
001822 => x"6163743A",
001823 => x"2073746E",
001824 => x"6F6C7469",
001825 => x"6E674067",
001826 => x"6F6F676C",
001827 => x"656D6169",
001828 => x"6C2E636F",
001829 => x"6D0D0A00",
001830 => x"28632920",
001831 => x"32303132",
001832 => x"20627920",
001833 => x"53746570",
001834 => x"68616E20",
001835 => x"4E6F6C74",
001836 => x"696E670D",
001837 => x"0A0D0A53",
001838 => x"656C6563",
001839 => x"743A2000",
001840 => x"0D0A0D0A",
001841 => x"5765276C",
001842 => x"6C207365",
001843 => x"6E642079",
001844 => x"6F752062",
001845 => x"61636B20",
001846 => x"2D20746F",
001847 => x"20746865",
001848 => x"20667574",
001849 => x"75726521",
001850 => x"2E0D0A0D",
001851 => x"0A000000",
001852 => x"202D2044",
001853 => x"6F63746F",
001854 => x"7220456D",
001855 => x"6D657420",
001856 => x"4C2E2042",
001857 => x"726F776E",
001858 => x"0D0A0D0A",
001859 => x"53656C65",
001860 => x"63743A20",
001861 => x"00000000",
001862 => x"20496E76",
001863 => x"616C6964",
001864 => x"206F7065",
001865 => x"72617469",
001866 => x"6F6E210D",
001867 => x"0A547279",
001868 => x"20616761",
001869 => x"696E3A20",
001870 => x"00000000",
001871 => x"0D0A0D0A",
001872 => x"2D3E2053",
001873 => x"74617274",
001874 => x"696E6720",
001875 => x"6170706C",
001876 => x"69636174",
001877 => x"696F6E2E",
001878 => x"2E2E0D0A",
001879 => x"0D0A0000",
001880 => x"0D0A0D0A",
001881 => x"41626F72",
001882 => x"74656421",
001883 => x"00000000",
others => x"F0013007"	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;