-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
	--bootloader sdram
000000 => x"EA000006",
000001 => x"EAFFFFFE",
000002 => x"EAFFFFFE",
000003 => x"EAFFFFFE",
000004 => x"EAFFFFFE",
000005 => x"E1A00000",
000006 => x"EAFFFFFE",
000007 => x"EAFFFFFE",
000008 => x"E59F0040",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA018",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"E1A04000",
000023 => x"E3A00000",
000024 => x"E1A0F004",
000025 => x"EAFFFFFE",
000026 => x"00002000",
000027 => x"0001084C",
000028 => x"E3E03A0F",
000029 => x"E5131FFB",
000030 => x"E20020FF",
000031 => x"E3A00001",
000032 => x"E0010210",
000033 => x"E1A0F00E",
000034 => x"E3E03A0F",
000035 => x"E5130FFB",
000036 => x"E1A0F00E",
000037 => x"E3E01A0F",
000038 => x"E5113FFF",
000039 => x"E20000FF",
000040 => x"E3A02001",
000041 => x"E1833012",
000042 => x"E5013FFF",
000043 => x"E1A0F00E",
000044 => x"E20000FF",
000045 => x"E3A02001",
000046 => x"E1A02012",
000047 => x"E3E01A0F",
000048 => x"E5113FFF",
000049 => x"E1E02002",
000050 => x"E0033002",
000051 => x"E5013FFF",
000052 => x"E1A0F00E",
000053 => x"E3E01A0F",
000054 => x"E5113FFF",
000055 => x"E20000FF",
000056 => x"E3A02001",
000057 => x"E0233012",
000058 => x"E5013FFF",
000059 => x"E1A0F00E",
000060 => x"E3E03A0F",
000061 => x"E5030FFF",
000062 => x"E1A0F00E",
000063 => x"E20000FF",
000064 => x"E3500007",
000065 => x"E92D4010",
000066 => x"E3A0C000",
000067 => x"E3E0E0FF",
000068 => x"E20110FF",
000069 => x"8A000011",
000070 => x"E2403004",
000071 => x"E20330FF",
000072 => x"E3500003",
000073 => x"E1A0E183",
000074 => x"E3E04A0F",
000075 => x"E1A0C180",
000076 => x"9A000007",
000077 => x"E3A030FF",
000078 => x"E1A03E13",
000079 => x"E5142F8B",
000080 => x"E1E03003",
000081 => x"E0022003",
000082 => x"E1822E11",
000083 => x"E5042F8B",
000084 => x"E8BD8010",
000085 => x"E3A030FF",
000086 => x"E1A03C13",
000087 => x"E1E0E003",
000088 => x"E3E02A0F",
000089 => x"E5123F8F",
000090 => x"E003300E",
000091 => x"E1833C11",
000092 => x"E5023F8F",
000093 => x"E8BD8010",
000094 => x"E20000FF",
000095 => x"E3500007",
000096 => x"E3A02000",
000097 => x"8A00000A",
000098 => x"E2403004",
000099 => x"E3500003",
000100 => x"E20320FF",
000101 => x"9A000005",
000102 => x"E3E03A0F",
000103 => x"E5130F8B",
000104 => x"E1A02182",
000105 => x"E1A00230",
000106 => x"E20000FF",
000107 => x"E1A0F00E",
000108 => x"E1A02180",
000109 => x"E3E03A0F",
000110 => x"E5130F8F",
000111 => x"E1A00230",
000112 => x"E20000FF",
000113 => x"E1A0F00E",
000114 => x"E3E02A0F",
000115 => x"E5123EFB",
000116 => x"E3130002",
000117 => x"E3E00000",
000118 => x"15120EFF",
000119 => x"E1A0F00E",
000120 => x"E3E02A0F",
000121 => x"E5123EFB",
000122 => x"E3130001",
000123 => x"0AFFFFFC",
000124 => x"E20030FF",
000125 => x"E5023EFF",
000126 => x"E1A0F00E",
000127 => x"E20000FF",
000128 => x"E3500001",
000129 => x"E3812B01",
000130 => x"03E03A0F",
000131 => x"E3811B09",
000132 => x"13E03A0F",
000133 => x"05031CFF",
000134 => x"15032CFF",
000135 => x"E1A0F00E",
000136 => x"E3E03A0F",
000137 => x"E5030CFB",
000138 => x"E1A0F00E",
000139 => x"E3E02A0F",
000140 => x"E5123CFF",
000141 => x"E3130C01",
000142 => x"1AFFFFFC",
000143 => x"E5020CEF",
000144 => x"E5123CFF",
000145 => x"E3833C01",
000146 => x"E5023CFF",
000147 => x"E3E02A0F",
000148 => x"E5123CFF",
000149 => x"E3130C01",
000150 => x"1AFFFFFC",
000151 => x"E5120CEF",
000152 => x"E1A0F00E",
000153 => x"E3E01A0F",
000154 => x"E5113CF7",
000155 => x"E20000FF",
000156 => x"E3A02001",
000157 => x"E1833012",
000158 => x"E5013CF7",
000159 => x"E1A0F00E",
000160 => x"E20000FF",
000161 => x"E3A02001",
000162 => x"E1A02012",
000163 => x"E3E01A0F",
000164 => x"E5113CF7",
000165 => x"E1E02002",
000166 => x"E0033002",
000167 => x"E5013CF7",
000168 => x"E1A0F00E",
000169 => x"E3E02A0F",
000170 => x"E5123BE7",
000171 => x"E1A01420",
000172 => x"E3C33080",
000173 => x"E5023BE7",
000174 => x"E5020BEF",
000175 => x"E5021BEB",
000176 => x"E5123BE7",
000177 => x"E3833080",
000178 => x"E5023BE7",
000179 => x"E1A0F00E",
000180 => x"E92D4030",
000181 => x"E3A0C090",
000182 => x"E20140FE",
000183 => x"E3E0EA0F",
000184 => x"E5DD500F",
000185 => x"E20000FF",
000186 => x"E50E4BE3",
000187 => x"E20110FF",
000188 => x"E50ECBFF",
000189 => x"E1A04002",
000190 => x"E203C0FF",
000191 => x"E51E3BFF",
000192 => x"E3130002",
000193 => x"1AFFFFFC",
000194 => x"E51E3BFF",
000195 => x"E3130080",
000196 => x"13E00000",
000197 => x"18BD8030",
000198 => x"E35C0000",
000199 => x"0A000012",
000200 => x"E24C3001",
000201 => x"E203C0FF",
000202 => x"E35C0001",
000203 => x"01A02424",
000204 => x"03E03A0F",
000205 => x"13E03A0F",
000206 => x"05032BE3",
000207 => x"15034BE3",
000208 => x"E3E02A0F",
000209 => x"E3A03010",
000210 => x"E5023BFF",
000211 => x"E5123BFF",
000212 => x"E3130002",
000213 => x"1AFFFFFC",
000214 => x"E5123BFF",
000215 => x"E3130080",
000216 => x"0AFFFFEC",
000217 => x"E3E00001",
000218 => x"E8BD8030",
000219 => x"E3500077",
000220 => x"1A00000C",
000221 => x"E3E03A0F",
000222 => x"E3A02050",
000223 => x"E5035BE3",
000224 => x"E5032BFF",
000225 => x"E1A02003",
000226 => x"E5123BFF",
000227 => x"E3130002",
000228 => x"1AFFFFFC",
000229 => x"E5123BFF",
000230 => x"E2130080",
000231 => x"08BD8030",
000232 => x"E3E00002",
000233 => x"E8BD8030",
000234 => x"E3500072",
000235 => x"13E00003",
000236 => x"18BD8030",
000237 => x"E3813001",
000238 => x"E3E02A0F",
000239 => x"E3A01090",
000240 => x"E5023BE3",
000241 => x"E5021BFF",
000242 => x"E5123BFF",
000243 => x"E3130002",
000244 => x"1AFFFFFC",
000245 => x"E5123BFF",
000246 => x"E3130080",
000247 => x"1AFFFFEF",
000248 => x"E3A03068",
000249 => x"E5023BFF",
000250 => x"E3E00A0F",
000251 => x"E5103BFF",
000252 => x"E3130002",
000253 => x"1AFFFFFC",
000254 => x"E5100BE3",
000255 => x"E8BD8030",
000256 => x"E20000FF",
000257 => x"E350000F",
000258 => x"979FF100",
000259 => x"EA00000F",
000260 => x"000104D0",
000261 => x"000104C8",
000262 => x"000104C0",
000263 => x"000104B8",
000264 => x"000104B0",
000265 => x"000104A8",
000266 => x"000104A0",
000267 => x"00010498",
000268 => x"00010490",
000269 => x"00010488",
000270 => x"00010480",
000271 => x"00010478",
000272 => x"00010470",
000273 => x"00010468",
000274 => x"00010460",
000275 => x"00010458",
000276 => x"E3A00000",
000277 => x"E1A0F00E",
000278 => x"EE1F0F1F",
000279 => x"E1A0F00E",
000280 => x"EE1E0F1E",
000281 => x"E1A0F00E",
000282 => x"EE1D0F1D",
000283 => x"E1A0F00E",
000284 => x"EE1C0F1C",
000285 => x"E1A0F00E",
000286 => x"EE1B0F1B",
000287 => x"E1A0F00E",
000288 => x"EE1A0F1A",
000289 => x"E1A0F00E",
000290 => x"EE190F19",
000291 => x"E1A0F00E",
000292 => x"EE180F18",
000293 => x"E1A0F00E",
000294 => x"EE170F17",
000295 => x"E1A0F00E",
000296 => x"EE160F16",
000297 => x"E1A0F00E",
000298 => x"EE150F15",
000299 => x"E1A0F00E",
000300 => x"EE140F14",
000301 => x"E1A0F00E",
000302 => x"EE130F13",
000303 => x"E1A0F00E",
000304 => x"EE120F12",
000305 => x"E1A0F00E",
000306 => x"EE110F11",
000307 => x"E1A0F00E",
000308 => x"EE100F10",
000309 => x"E1A0F00E",
000310 => x"E20110FF",
000311 => x"E2411006",
000312 => x"E3510007",
000313 => x"979FF101",
000314 => x"EA000008",
000315 => x"00010514",
000316 => x"00010510",
000317 => x"00010510",
000318 => x"00010510",
000319 => x"00010510",
000320 => x"0001051C",
000321 => x"00010524",
000322 => x"0001050C",
000323 => x"EE0D0F1D",
000324 => x"E1A0F00E",
000325 => x"EE060F16",
000326 => x"E1A0F00E",
000327 => x"EE0B0F1B",
000328 => x"E1A0F00E",
000329 => x"EE0C0F1C",
000330 => x"E1A0F00E",
000331 => x"E92D4010",
000332 => x"E1A04000",
000333 => x"E5D00000",
000334 => x"E3500000",
000335 => x"1A000003",
000336 => x"EA000005",
000337 => x"E5F40001",
000338 => x"E3500000",
000339 => x"0A000002",
000340 => x"EBFFFF22",
000341 => x"E3500000",
000342 => x"CAFFFFF9",
000343 => x"E1A00004",
000344 => x"E8BD8010",
000345 => x"E92D4070",
000346 => x"E2514000",
000347 => x"E1A05000",
000348 => x"E20260FF",
000349 => x"DA00000B",
000350 => x"EBFFFF12",
000351 => x"E3700001",
000352 => x"E20030FF",
000353 => x"0A000005",
000354 => x"E3560001",
000355 => x"E5C53000",
000356 => x"E1A00003",
000357 => x"E2855001",
000358 => x"0A000005",
000359 => x"E2444001",
000360 => x"E3540000",
000361 => x"CAFFFFF3",
000362 => x"E59F300C",
000363 => x"E5C53000",
000364 => x"E8BD8070",
000365 => x"EBFFFF09",
000366 => x"EAFFFFF7",
000367 => x"00011188",
000368 => x"E92D4030",
000369 => x"E2514000",
000370 => x"E1A05000",
000371 => x"D8BD8030",
000372 => x"E4D50001",
000373 => x"EBFFFF01",
000374 => x"E2544001",
000375 => x"1AFFFFFB",
000376 => x"E8BD8030",
000377 => x"E92D4010",
000378 => x"E20240FF",
000379 => x"E3540008",
000380 => x"83A04008",
000381 => x"8A000001",
000382 => x"E3540000",
000383 => x"03A04001",
000384 => x"E1A02001",
000385 => x"E1A0E004",
000386 => x"E1A0310E",
000387 => x"E35E0001",
000388 => x"E2433004",
000389 => x"E1A0C000",
000390 => x"81A0C330",
000391 => x"E24E3001",
000392 => x"E20CC00F",
000393 => x"E203E0FF",
000394 => x"E35C0009",
000395 => x"E28C3030",
000396 => x"828C3037",
000397 => x"E35E0000",
000398 => x"E4C23001",
000399 => x"1AFFFFF1",
000400 => x"E2443001",
000401 => x"E20330FF",
000402 => x"E0813003",
000403 => x"E5C3E001",
000404 => x"E8BD8010",
000405 => x"E92D4010",
000406 => x"E1A04000",
000407 => x"E3540007",
000408 => x"E3A01010",
000409 => x"E3A00001",
000410 => x"9A000001",
000411 => x"E3A00000",
000412 => x"E8BD8010",
000413 => x"EBFFFEE0",
000414 => x"E3A00006",
000415 => x"EBFFFEF8",
000416 => x"E3A00000",
000417 => x"EBFFFEE8",
000418 => x"E1A00584",
000419 => x"E8BD4010",
000420 => x"EAFFFEE5",
000421 => x"E0603280",
000422 => x"E0800103",
000423 => x"E0800100",
000424 => x"E1A00200",
000425 => x"E3500000",
000426 => x"D1A0F00E",
000427 => x"E1A00000",
000428 => x"E2500001",
000429 => x"1AFFFFFC",
000430 => x"E1A0F00E",
000431 => x"E212C0FF",
000432 => x"0A00000B",
000433 => x"E5D02000",
000434 => x"E5D13000",
000435 => x"E1520003",
000436 => x"0A000004",
000437 => x"EA000008",
000438 => x"E5F02001",
000439 => x"E5F13001",
000440 => x"E1520003",
000441 => x"1A000004",
000442 => x"E24C3001",
000443 => x"E213C0FF",
000444 => x"1AFFFFF8",
000445 => x"E3A00001",
000446 => x"E1A0F00E",
000447 => x"E3A00000",
000448 => x"E1A0F00E",
000449 => x"E92D4030",
000450 => x"E1A04081",
000451 => x"E3540000",
000452 => x"E1A05000",
000453 => x"D3A00000",
000454 => x"D8BD8030",
000455 => x"E3A00000",
000456 => x"E1A01000",
000457 => x"E7D12005",
000458 => x"E2423030",
000459 => x"E082C200",
000460 => x"E3530009",
000461 => x"E242E041",
000462 => x"924C0030",
000463 => x"9A000007",
000464 => x"E0823200",
000465 => x"E35E0005",
000466 => x"E242C061",
000467 => x"92430037",
000468 => x"9A000002",
000469 => x"E0823200",
000470 => x"E35C0005",
000471 => x"92430057",
000472 => x"E2811001",
000473 => x"E1510004",
000474 => x"1AFFFFED",
000475 => x"E8BD8030",
000476 => x"E52DE004",
000477 => x"E59F0074",
000478 => x"EBFFFF6B",
000479 => x"E59F0070",
000480 => x"EBFFFF69",
000481 => x"E59F006C",
000482 => x"EBFFFF67",
000483 => x"E59F0068",
000484 => x"EBFFFF65",
000485 => x"E59F0064",
000486 => x"EBFFFF63",
000487 => x"E59F0060",
000488 => x"EBFFFF61",
000489 => x"E59F005C",
000490 => x"EBFFFF5F",
000491 => x"E59F0058",
000492 => x"EBFFFF5D",
000493 => x"E59F0054",
000494 => x"EBFFFF5B",
000495 => x"E59F0050",
000496 => x"EBFFFF59",
000497 => x"E59F004C",
000498 => x"EBFFFF57",
000499 => x"E59F0048",
000500 => x"EBFFFF55",
000501 => x"E59F0044",
000502 => x"EBFFFF53",
000503 => x"E59F0040",
000504 => x"EBFFFF51",
000505 => x"E59F003C",
000506 => x"E49DE004",
000507 => x"EAFFFF4E",
000508 => x"0001118C",
000509 => x"000111D8",
000510 => x"00011220",
000511 => x"00011268",
000512 => x"000112B0",
000513 => x"000112F8",
000514 => x"00011340",
000515 => x"00011380",
000516 => x"000113B8",
000517 => x"000113DC",
000518 => x"00011424",
000519 => x"00011490",
000520 => x"000114C8",
000521 => x"0001152C",
000522 => x"00011590",
000523 => x"E5D03003",
000524 => x"E5D02002",
000525 => x"E5D01000",
000526 => x"E1833402",
000527 => x"E5D00001",
000528 => x"E1833C01",
000529 => x"E1830800",
000530 => x"E1A0F00E",
000531 => x"E92D47F0",
000532 => x"E3A00000",
000533 => x"E24DD018",
000534 => x"EBFFFE24",
000535 => x"E3A0100D",
000536 => x"E3A000C3",
000537 => x"EBFFFF1B",
000538 => x"E3A00063",
000539 => x"EBFFFE8C",
000540 => x"E3A00006",
000541 => x"EBFFFEE1",
000542 => x"E3A01006",
000543 => x"E3800008",
000544 => x"EBFFFF14",
000545 => x"E3A0000D",
000546 => x"EBFFFEDC",
000547 => x"E1A008A0",
000548 => x"E1E00000",
000549 => x"E200000F",
000550 => x"E3500001",
000551 => x"03A04030",
000552 => x"028DA006",
000553 => x"028D900F",
000554 => x"0A00001A",
000555 => x"E3500002",
000556 => x"0A000077",
000557 => x"EBFFFFAD",
000558 => x"E28DA006",
000559 => x"E59F0808",
000560 => x"EBFFFF19",
000561 => x"E1A0100A",
000562 => x"E3A02008",
000563 => x"E28D0014",
000564 => x"EBFFFF43",
000565 => x"E1A0000A",
000566 => x"EBFFFF13",
000567 => x"E59F07EC",
000568 => x"EBFFFF11",
000569 => x"E59F07E8",
000570 => x"EBFFFF0F",
000571 => x"E1A0100A",
000572 => x"E3A02008",
000573 => x"E3A00301",
000574 => x"EBFFFF39",
000575 => x"E1A0000A",
000576 => x"EBFFFF09",
000577 => x"E59F07C4",
000578 => x"EBFFFF07",
000579 => x"E28D900F",
000580 => x"EBFFFE2C",
000581 => x"E1A04000",
000582 => x"E3A0000D",
000583 => x"EBFFFEB7",
000584 => x"E3100801",
000585 => x"03A06001",
000586 => x"03A040A0",
000587 => x"1A00003C",
000588 => x"E3A05000",
000589 => x"E59F079C",
000590 => x"EBFFFEFB",
000591 => x"E1A01004",
000592 => x"E1A02005",
000593 => x"E3A03002",
000594 => x"E3A00072",
000595 => x"E58D5000",
000596 => x"EBFFFE5E",
000597 => x"E1A01004",
000598 => x"E5CD000F",
000599 => x"E3A02001",
000600 => x"E3A03002",
000601 => x"E3A00072",
000602 => x"E58D5000",
000603 => x"EBFFFE57",
000604 => x"E3A02002",
000605 => x"E1A03002",
000606 => x"E5CD0010",
000607 => x"E1A01004",
000608 => x"E3A00072",
000609 => x"E58D5000",
000610 => x"EBFFFE50",
000611 => x"E3A03002",
000612 => x"E5CD0011",
000613 => x"E1A01004",
000614 => x"E3A00072",
000615 => x"E3A02003",
000616 => x"E58D5000",
000617 => x"EBFFFE49",
000618 => x"E5DD300F",
000619 => x"E20000FF",
000620 => x"E3530053",
000621 => x"E5CD0012",
000622 => x"1A000002",
000623 => x"E5DD3010",
000624 => x"E353004D",
000625 => x"0A00006A",
000626 => x"E59F070C",
000627 => x"EBFFFED6",
000628 => x"E3560000",
000629 => x"0AFFFFCD",
000630 => x"E59F0700",
000631 => x"EBFFFED2",
000632 => x"E3A0100D",
000633 => x"E3A00000",
000634 => x"EBFFFEBA",
000635 => x"E59F06F0",
000636 => x"EBFFFECD",
000637 => x"E3A00006",
000638 => x"EBFFFE80",
000639 => x"E3A01006",
000640 => x"E3C00008",
000641 => x"EBFFFEB3",
000642 => x"E59F06D8",
000643 => x"EBFFFEC6",
000644 => x"E3A00301",
000645 => x"EBFFFD8F",
000646 => x"E59F06CC",
000647 => x"EBFFFEC2",
000648 => x"EAFFFFFE",
000649 => x"E3540034",
000650 => x"0A000029",
000651 => x"CA00001C",
000652 => x"E3540031",
000653 => x"0A000036",
000654 => x"DA00009B",
000655 => x"E3540032",
000656 => x"0A0000A5",
000657 => x"E3540033",
000658 => x"1A00009B",
000659 => x"E1A00004",
000660 => x"EBFFFDE2",
000661 => x"E59F0694",
000662 => x"EBFFFEB3",
000663 => x"E1A00009",
000664 => x"E3A01002",
000665 => x"E3A02001",
000666 => x"EBFFFEBD",
000667 => x"E3A01002",
000668 => x"E1A00009",
000669 => x"EBFFFF22",
000670 => x"E21010FF",
000671 => x"11A04001",
000672 => x"13A06000",
000673 => x"1AFFFFA9",
000674 => x"E59F0664",
000675 => x"EBFFFEA6",
000676 => x"EAFFFF9E",
000677 => x"E3A04033",
000678 => x"E28DA006",
000679 => x"E28D900F",
000680 => x"EAFFFF9C",
000681 => x"E3540066",
000682 => x"0A00002A",
000683 => x"DA0000B0",
000684 => x"E3540068",
000685 => x"0A000112",
000686 => x"E3540072",
000687 => x"1A00007E",
000688 => x"E1A00004",
000689 => x"EBFFFDC5",
000690 => x"E3A006FF",
000691 => x"E280F20F",
000692 => x"EAFFFFFE",
000693 => x"E1A00004",
000694 => x"EBFFFDC0",
000695 => x"E59F060C",
000696 => x"EBFFFE91",
000697 => x"E1A00009",
000698 => x"E3A01002",
000699 => x"E3A02001",
000700 => x"EBFFFE9B",
000701 => x"E1A00009",
000702 => x"E3A01002",
000703 => x"EBFFFF00",
000704 => x"E21080FF",
000705 => x"1A0000A7",
000706 => x"E59F05E8",
000707 => x"EBFFFE86",
000708 => x"EAFFFF7E",
000709 => x"E1A00004",
000710 => x"EBFFFDB0",
000711 => x"E59F05D8",
000712 => x"EBFFFE81",
000713 => x"E1A00009",
000714 => x"E3A01004",
000715 => x"E3A02000",
000716 => x"EBFFFE8B",
000717 => x"E5DD300F",
000718 => x"E3530053",
000719 => x"1A000002",
000720 => x"E5DD3010",
000721 => x"E353004D",
000722 => x"0A0000F1",
000723 => x"E59F05AC",
000724 => x"EBFFFE75",
000725 => x"EAFFFF6D",
000726 => x"E1A00004",
000727 => x"EBFFFD9F",
000728 => x"E59F059C",
000729 => x"EBFFFE70",
000730 => x"E59F0598",
000731 => x"EBFFFE6E",
000732 => x"EAFFFF66",
000733 => x"E5DD3011",
000734 => x"E3530042",
000735 => x"1AFFFF91",
000736 => x"E3500052",
000737 => x"1AFFFF8F",
000738 => x"E1A01004",
000739 => x"E3A02004",
000740 => x"E2433040",
000741 => x"E2800020",
000742 => x"E58D5000",
000743 => x"EBFFFDCB",
000744 => x"E1A01004",
000745 => x"E5CD000F",
000746 => x"E3A02005",
000747 => x"E3A03002",
000748 => x"E3A00072",
000749 => x"E58D5000",
000750 => x"EBFFFDC4",
000751 => x"E1A01004",
000752 => x"E5CD0010",
000753 => x"E3A02006",
000754 => x"E3A03002",
000755 => x"E3A00072",
000756 => x"E58D5000",
000757 => x"EBFFFDBD",
000758 => x"E1A01004",
000759 => x"E5CD0011",
000760 => x"E3A02007",
000761 => x"E3A03002",
000762 => x"E3A00072",
000763 => x"E58D5000",
000764 => x"EBFFFDB6",
000765 => x"E5CD0012",
000766 => x"E1A00009",
000767 => x"EBFFFF0A",
000768 => x"E3700004",
000769 => x"E58D0014",
000770 => x"0A000024",
000771 => x"E1A06005",
000772 => x"E2852008",
000773 => x"E1A01004",
000774 => x"E3A03002",
000775 => x"E3A00072",
000776 => x"E58D6000",
000777 => x"EBFFFDA9",
000778 => x"E2852009",
000779 => x"E5CD000F",
000780 => x"E1A01004",
000781 => x"E3A03002",
000782 => x"E3A00072",
000783 => x"E58D6000",
000784 => x"EBFFFDA2",
000785 => x"E285200A",
000786 => x"E5CD0010",
000787 => x"E1A01004",
000788 => x"E3A03002",
000789 => x"E3A00072",
000790 => x"E58D6000",
000791 => x"EBFFFD9B",
000792 => x"E285200B",
000793 => x"E3A03002",
000794 => x"E5CD0011",
000795 => x"E1A01004",
000796 => x"E3A00072",
000797 => x"E58D6000",
000798 => x"EBFFFD94",
000799 => x"E5CD0012",
000800 => x"E1A00009",
000801 => x"EBFFFEE8",
000802 => x"E4850004",
000803 => x"E59D3014",
000804 => x"E2833004",
000805 => x"E1530005",
000806 => x"13550902",
000807 => x"3AFFFFDB",
000808 => x"E59F0464",
000809 => x"EBFFFE20",
000810 => x"EAFFFF4A",
000811 => x"E3740001",
000812 => x"0AFFFF16",
000813 => x"E3540030",
000814 => x"0A000004",
000815 => x"E20400FF",
000816 => x"EBFFFD46",
000817 => x"E59F0444",
000818 => x"EBFFFE17",
000819 => x"EAFFFF0F",
000820 => x"E1A00004",
000821 => x"EBFFFD41",
000822 => x"EAFFFF3E",
000823 => x"E1A00004",
000824 => x"EBFFFD3E",
000825 => x"E59F0428",
000826 => x"EBFFFE0F",
000827 => x"EBFFFD35",
000828 => x"E3700001",
000829 => x"0AFFFFFC",
000830 => x"EBFFFD32",
000831 => x"E3700001",
000832 => x"1AFFFFFC",
000833 => x"E3A05301",
000834 => x"E5950000",
000835 => x"E1A0100A",
000836 => x"E3A02008",
000837 => x"EBFFFE32",
000838 => x"E5DD0006",
000839 => x"E3500000",
000840 => x"0A000005",
000841 => x"E3A04000",
000842 => x"E2844001",
000843 => x"EBFFFD2B",
000844 => x"E7D4000A",
000845 => x"E3500000",
000846 => x"1AFFFFFA",
000847 => x"E3A00020",
000848 => x"EBFFFD26",
000849 => x"EBFFFD1F",
000850 => x"E3700001",
000851 => x"1A000005",
000852 => x"E3A03301",
000853 => x"E2833E9E",
000854 => x"E2855004",
000855 => x"E2833004",
000856 => x"E1550003",
000857 => x"1AFFFFE7",
000858 => x"E59F03A8",
000859 => x"EBFFFDEE",
000860 => x"EAFFFEE6",
000861 => x"E3540035",
000862 => x"0A00009C",
000863 => x"E3540061",
000864 => x"1AFFFFCD",
000865 => x"E1A00004",
000866 => x"EBFFFD14",
000867 => x"E59F0388",
000868 => x"EBFFFDE5",
000869 => x"E59F0384",
000870 => x"EBFFFDE3",
000871 => x"E59F0380",
000872 => x"EBFFFDE1",
000873 => x"EAFFFED9",
000874 => x"E59F0378",
000875 => x"EBFFFDDE",
000876 => x"E1A00009",
000877 => x"E3A01004",
000878 => x"E3A02000",
000879 => x"EBFFFDE8",
000880 => x"E5DD300F",
000881 => x"E3530053",
000882 => x"1A000002",
000883 => x"E5DD2010",
000884 => x"E352004D",
000885 => x"0A000004",
000886 => x"E59F034C",
000887 => x"EBFFFDD2",
000888 => x"E59F0348",
000889 => x"EBFFFDD0",
000890 => x"EAFFFEC8",
000891 => x"E5DD1011",
000892 => x"E3510042",
000893 => x"1AFFFFF7",
000894 => x"E5DD0012",
000895 => x"E3500052",
000896 => x"1AFFFFF4",
000897 => x"E3A04000",
000898 => x"E5C43000",
000899 => x"E1A00000",
000900 => x"E5C42001",
000901 => x"E1A00000",
000902 => x"E5C41002",
000903 => x"E1A00000",
000904 => x"E5C40003",
000905 => x"E1A00000",
000906 => x"E241103E",
000907 => x"E1A00009",
000908 => x"E1A02004",
000909 => x"EBFFFDCA",
000910 => x"E5DD300F",
000911 => x"E5C43004",
000912 => x"E5DD2010",
000913 => x"E5C42005",
000914 => x"E5DD3011",
000915 => x"E5C43006",
000916 => x"E5DD2012",
000917 => x"E1A00009",
000918 => x"E5C42007",
000919 => x"EBFFFE72",
000920 => x"E3A03CFF",
000921 => x"E28330FC",
000922 => x"E1500003",
000923 => x"E1A05000",
000924 => x"8A00008B",
000925 => x"E3700004",
000926 => x"12844008",
000927 => x"1280600B",
000928 => x"0A000006",
000929 => x"EBFFFCCF",
000930 => x"E3700001",
000931 => x"0AFFFFFC",
000932 => x"E1560004",
000933 => x"E5C40000",
000934 => x"E2844001",
000935 => x"1AFFFFF8",
000936 => x"E59F028C",
000937 => x"EBFFFDA0",
000938 => x"E59F0288",
000939 => x"EBFFFD9E",
000940 => x"E375000C",
000941 => x"0A00000F",
000942 => x"E3A04000",
000943 => x"E285700C",
000944 => x"E1A06004",
000945 => x"E5D45000",
000946 => x"E3A00077",
000947 => x"E1A01008",
000948 => x"E1A02006",
000949 => x"E3A03002",
000950 => x"E58D5000",
000951 => x"EBFFFCFB",
000952 => x"E3500000",
000953 => x"1AFFFFF7",
000954 => x"E2844001",
000955 => x"E1570004",
000956 => x"E1A06004",
000957 => x"1AFFFFF2",
000958 => x"E59F023C",
000959 => x"EBFFFD8A",
000960 => x"EAFFFFB6",
000961 => x"E1A00004",
000962 => x"EBFFFCB4",
000963 => x"EBFFFE17",
000964 => x"EAFFFE7E",
000965 => x"E5DD3011",
000966 => x"E3530042",
000967 => x"1AFFFF0A",
000968 => x"E5DD3012",
000969 => x"E3530052",
000970 => x"1AFFFF07",
000971 => x"E3A01004",
000972 => x"E3A02000",
000973 => x"E1A00009",
000974 => x"EBFFFD89",
000975 => x"E1A00009",
000976 => x"EBFFFE39",
000977 => x"E3A03402",
000978 => x"E2433008",
000979 => x"E1500003",
000980 => x"E58D0014",
000981 => x"8A00004F",
000982 => x"E2804301",
000983 => x"E2844004",
000984 => x"E3540301",
000985 => x"0A00000A",
000986 => x"E3A05301",
000987 => x"E3A01004",
000988 => x"E3A02000",
000989 => x"E1A00009",
000990 => x"EBFFFD79",
000991 => x"E1A00009",
000992 => x"EBFFFE29",
000993 => x"E4850004",
000994 => x"E1550004",
000995 => x"1AFFFFF6",
000996 => x"E1A04005",
000997 => x"E59F01A4",
000998 => x"EBFFFD63",
000999 => x"E1A0100A",
001000 => x"E3A02008",
001001 => x"E1A00004",
001002 => x"EBFFFD8D",
001003 => x"E1A0000A",
001004 => x"EBFFFD5D",
001005 => x"E59F0188",
001006 => x"EBFFFD5B",
001007 => x"E59F0184",
001008 => x"EBFFFD59",
001009 => x"E59F0180",
001010 => x"EBFFFD57",
001011 => x"E1A00004",
001012 => x"E1A0100A",
001013 => x"E3A02008",
001014 => x"EBFFFD81",
001015 => x"E1A0000A",
001016 => x"EBFFFD51",
001017 => x"E59F0158",
001018 => x"EBFFFD4F",
001019 => x"EAFFFE47",
001020 => x"E1A00004",
001021 => x"EBFFFC79",
001022 => x"E59F0150",
001023 => x"EBFFFD4A",
001024 => x"E1A00009",
001025 => x"E3A01002",
001026 => x"E3A02001",
001027 => x"EBFFFD54",
001028 => x"E1A00009",
001029 => x"E3A01002",
001030 => x"EBFFFDB9",
001031 => x"E21060FF",
001032 => x"0AFFFE98",
001033 => x"E59F0128",
001034 => x"EBFFFD3F",
001035 => x"E59F0124",
001036 => x"EBFFFD3D",
001037 => x"EBFFFC63",
001038 => x"E3700001",
001039 => x"0AFFFFFC",
001040 => x"EBFFFC60",
001041 => x"E3700001",
001042 => x"1AFFFFFC",
001043 => x"E3A05000",
001044 => x"EA000001",
001045 => x"E3540000",
001046 => x"AA000014",
001047 => x"E3A0C000",
001048 => x"E1A02005",
001049 => x"E1A01006",
001050 => x"E3A03002",
001051 => x"E3A00072",
001052 => x"E58DC000",
001053 => x"EBFFFC95",
001054 => x"E1A04000",
001055 => x"EBFFFC51",
001056 => x"E3700001",
001057 => x"E1A00004",
001058 => x"0AFFFFF1",
001059 => x"E59F00C8",
001060 => x"EBFFFD25",
001061 => x"EAFFFF33",
001062 => x"E59F00C0",
001063 => x"EBFFFD22",
001064 => x"EAFFFE1A",
001065 => x"E59F00B8",
001066 => x"EBFFFD1F",
001067 => x"EAFFFE17",
001068 => x"EBFFFC4A",
001069 => x"E3A03801",
001070 => x"E2855001",
001071 => x"E2433001",
001072 => x"E1550003",
001073 => x"1AFFFFE4",
001074 => x"EAFFFF26",
001075 => x"000115E0",
001076 => x"000115F8",
001077 => x"00011600",
001078 => x"000117D4",
001079 => x"00011838",
001080 => x"00011B98",
001081 => x"00011BBC",
001082 => x"00011BEC",
001083 => x"00011C10",
001084 => x"00011778",
001085 => x"000117B4",
001086 => x"00011864",
001087 => x"00011610",
001088 => x"000116E4",
001089 => x"00011B1C",
001090 => x"00011B4C",
001091 => x"00011824",
001092 => x"00011B74",
001093 => x"0001170C",
001094 => x"00011754",
001095 => x"00011A38",
001096 => x"00011A6C",
001097 => x"00011AD8",
001098 => x"00011884",
001099 => x"00011950",
001100 => x"00011B68",
001101 => x"00011908",
001102 => x"00011920",
001103 => x"00011940",
001104 => x"000116AC",
001105 => x"000116C0",
001106 => x"000116C4",
001107 => x"000116D4",
001108 => x"00011974",
001109 => x"000119B0",
001110 => x"000119F0",
001111 => x"00011C2C",
001112 => x"00011684",
001113 => x"000118E4",
001114 => x"E10F3000",
001115 => x"E3C330C0",
001116 => x"E129F003",
001117 => x"E1A0F00E",
001118 => x"E10F3000",
001119 => x"E38330C0",
001120 => x"E129F003",
001121 => x"E1A0F00E",
001122 => x"00000000",
001123 => x"0D0A0D0A",
001124 => x"0D0A2B2D",
001125 => x"2D2D2D2D",
001126 => x"2D2D2D2D",
001127 => x"2D2D2D2D",
001128 => x"2D2D2D2D",
001129 => x"2D2D2D2D",
001130 => x"2D2D2D2D",
001131 => x"2D2D2D2D",
001132 => x"2D2D2D2D",
001133 => x"2D2D2D2D",
001134 => x"2D2D2D2D",
001135 => x"2D2D2D2D",
001136 => x"2D2D2D2D",
001137 => x"2D2D2D2D",
001138 => x"2D2D2D2D",
001139 => x"2D2D2D2D",
001140 => x"2D2D2D2B",
001141 => x"0D0A0000",
001142 => x"7C202020",
001143 => x"203C3C3C",
001144 => x"2053544F",
001145 => x"524D2043",
001146 => x"6F726520",
001147 => x"50726F63",
001148 => x"6573736F",
001149 => x"72205379",
001150 => x"7374656D",
001151 => x"202D2042",
001152 => x"79205374",
001153 => x"65706861",
001154 => x"6E204E6F",
001155 => x"6C74696E",
001156 => x"67203E3E",
001157 => x"3E202020",
001158 => x"207C0D0A",
001159 => x"00000000",
001160 => x"2B2D2D2D",
001161 => x"2D2D2D2D",
001162 => x"2D2D2D2D",
001163 => x"2D2D2D2D",
001164 => x"2D2D2D2D",
001165 => x"2D2D2D2D",
001166 => x"2D2D2D2D",
001167 => x"2D2D2D2D",
001168 => x"2D2D2D2D",
001169 => x"2D2D2D2D",
001170 => x"2D2D2D2D",
001171 => x"2D2D2D2D",
001172 => x"2D2D2D2D",
001173 => x"2D2D2D2D",
001174 => x"2D2D2D2D",
001175 => x"2D2D2D2D",
001176 => x"2D2B0D0A",
001177 => x"00000000",
001178 => x"7C202020",
001179 => x"20202020",
001180 => x"2020426F",
001181 => x"6F746C6F",
001182 => x"61646572",
001183 => x"20666F72",
001184 => x"2053544F",
001185 => x"524D2053",
001186 => x"6F432020",
001187 => x"20566572",
001188 => x"73696F6E",
001189 => x"3A203230",
001190 => x"31323035",
001191 => x"32342D44",
001192 => x"20202020",
001193 => x"20202020",
001194 => x"207C0D0A",
001195 => x"00000000",
001196 => x"7C202020",
001197 => x"20202020",
001198 => x"20202020",
001199 => x"20202020",
001200 => x"436F6E74",
001201 => x"6163743A",
001202 => x"2073746E",
001203 => x"6F6C7469",
001204 => x"6E674067",
001205 => x"6F6F676C",
001206 => x"656D6169",
001207 => x"6C2E636F",
001208 => x"6D202020",
001209 => x"20202020",
001210 => x"20202020",
001211 => x"20202020",
001212 => x"207C0D0A",
001213 => x"00000000",
001214 => x"2B2D2D2D",
001215 => x"2D2D2D2D",
001216 => x"2D2D2D2D",
001217 => x"2D2D2D2D",
001218 => x"2D2D2D2D",
001219 => x"2D2D2D2D",
001220 => x"2D2D2D2D",
001221 => x"2D2D2D2D",
001222 => x"2D2D2D2D",
001223 => x"2D2D2D2D",
001224 => x"2D2D2D2D",
001225 => x"2D2D2D2D",
001226 => x"2D2D2D2D",
001227 => x"2D2D2D2D",
001228 => x"2D2D2D2D",
001229 => x"2D2D2D2D",
001230 => x"2D2B0D0A",
001231 => x"0D0A0000",
001232 => x"636F6E6E",
001233 => x"65637465",
001234 => x"6420746F",
001235 => x"20493243",
001236 => x"5F434F4E",
001237 => x"54524F4C",
001238 => x"4C45525F",
001239 => x"302C206F",
001240 => x"70657261",
001241 => x"74696E67",
001242 => x"20667265",
001243 => x"7175656E",
001244 => x"63792069",
001245 => x"73203130",
001246 => x"306B487A",
001247 => x"2C0D0A00",
001248 => x"6D617869",
001249 => x"6D756D20",
001250 => x"45455052",
001251 => x"4F4D2073",
001252 => x"697A6520",
001253 => x"3D203635",
001254 => x"35333620",
001255 => x"62797465",
001256 => x"203D3E20",
001257 => x"31362062",
001258 => x"69742061",
001259 => x"64647265",
001260 => x"73736573",
001261 => x"2C0D0A00",
001262 => x"66697865",
001263 => x"6420626F",
001264 => x"6F742064",
001265 => x"65766963",
001266 => x"65206164",
001267 => x"64726573",
001268 => x"733A2030",
001269 => x"7841300D",
001270 => x"0A0D0A00",
001271 => x"426F6F74",
001272 => x"20454550",
001273 => x"524F4D3A",
001274 => x"20323478",
001275 => x"786E6E6E",
001276 => x"20286C69",
001277 => x"6B652032",
001278 => x"34414136",
001279 => x"34292C20",
001280 => x"37206269",
001281 => x"74206164",
001282 => x"64726573",
001283 => x"73202B20",
001284 => x"646F6E74",
001285 => x"2D636172",
001286 => x"65206269",
001287 => x"742C0D0A",
001288 => x"00000000",
001289 => x"203C2057",
001290 => x"656C636F",
001291 => x"6D652074",
001292 => x"6F207468",
001293 => x"65205354",
001294 => x"4F524D20",
001295 => x"536F4320",
001296 => x"626F6F74",
001297 => x"6C6F6164",
001298 => x"65722063",
001299 => x"6F6E736F",
001300 => x"6C652120",
001301 => x"3E0D0A20",
001302 => x"3C205365",
001303 => x"6C656374",
001304 => x"20616E20",
001305 => x"6F706572",
001306 => x"6174696F",
001307 => x"6E206672",
001308 => x"6F6D2074",
001309 => x"6865206D",
001310 => x"656E7520",
001311 => x"62656C6F",
001312 => x"77206F72",
001313 => x"20707265",
001314 => x"7373203E",
001315 => x"0D0A0000",
001316 => x"203C2074",
001317 => x"68652062",
001318 => x"6F6F7420",
001319 => x"6B657920",
001320 => x"666F7220",
001321 => x"696D6D65",
001322 => x"64696174",
001323 => x"65206170",
001324 => x"706C6963",
001325 => x"6174696F",
001326 => x"6E207374",
001327 => x"6172742E",
001328 => x"203E0D0A",
001329 => x"0D0A0000",
001330 => x"2030202D",
001331 => x"20626F6F",
001332 => x"74206672",
001333 => x"6F6D2063",
001334 => x"6F726520",
001335 => x"52414D20",
001336 => x"28737461",
001337 => x"72742061",
001338 => x"70706C69",
001339 => x"63617469",
001340 => x"6F6E290D",
001341 => x"0A203120",
001342 => x"2D207072",
001343 => x"6F677261",
001344 => x"6D20636F",
001345 => x"72652052",
001346 => x"414D2076",
001347 => x"69612055",
001348 => x"4152545F",
001349 => x"300D0A20",
001350 => x"32202D20",
001351 => x"636F7265",
001352 => x"2052414D",
001353 => x"2064756D",
001354 => x"700D0A00",
001355 => x"2033202D",
001356 => x"20626F6F",
001357 => x"74206672",
001358 => x"6F6D2049",
001359 => x"32432045",
001360 => x"4550524F",
001361 => x"4D0D0A20",
001362 => x"34202D20",
001363 => x"70726F67",
001364 => x"72616D20",
001365 => x"49324320",
001366 => x"45455052",
001367 => x"4F4D2076",
001368 => x"69612055",
001369 => x"4152545F",
001370 => x"300D0A20",
001371 => x"35202D20",
001372 => x"73686F77",
001373 => x"20636F6E",
001374 => x"74656E74",
001375 => x"206F6620",
001376 => x"49324320",
001377 => x"45455052",
001378 => x"4F4D0D0A",
001379 => x"00000000",
001380 => x"2061202D",
001381 => x"20617574",
001382 => x"6F6D6174",
001383 => x"69632062",
001384 => x"6F6F7420",
001385 => x"636F6E66",
001386 => x"69677572",
001387 => x"6174696F",
001388 => x"6E0D0A20",
001389 => x"68202D20",
001390 => x"68656C70",
001391 => x"0D0A2072",
001392 => x"202D2072",
001393 => x"65737461",
001394 => x"72742073",
001395 => x"79737465",
001396 => x"6D0D0A0D",
001397 => x"0A53656C",
001398 => x"6563743A",
001399 => x"20000000",
001400 => x"41646472",
001401 => x"65737320",
001402 => x"6F662061",
001403 => x"64725F62",
001404 => x"75666665",
001405 => x"723A2000",
001406 => x"200A0D20",
001407 => x"00000000",
001408 => x"204C6F61",
001409 => x"64204164",
001410 => x"64726573",
001411 => x"733A2000",
001412 => x"0D0A0D0A",
001413 => x"4170706C",
001414 => x"69636174",
001415 => x"696F6E20",
001416 => x"77696C6C",
001417 => x"20737461",
001418 => x"72742061",
001419 => x"75746F6D",
001420 => x"61746963",
001421 => x"616C6C79",
001422 => x"20616674",
001423 => x"65722064",
001424 => x"6F776E6C",
001425 => x"6F61642E",
001426 => x"0D0A2D3E",
001427 => x"20576169",
001428 => x"74696E67",
001429 => x"20666F72",
001430 => x"20277374",
001431 => x"6F726D5F",
001432 => x"70726F67",
001433 => x"72616D2E",
001434 => x"62696E27",
001435 => x"20696E20",
001436 => x"62797465",
001437 => x"2D737472",
001438 => x"65616D20",
001439 => x"6D6F6465",
001440 => x"2E2E2E00",
001441 => x"20534452",
001442 => x"414D2045",
001443 => x"52524F52",
001444 => x"21205072",
001445 => x"6F677261",
001446 => x"6D206669",
001447 => x"6C652074",
001448 => x"6F6F2062",
001449 => x"6967210D",
001450 => x"0A0D0A00",
001451 => x"4C617374",
001452 => x"206D656D",
001453 => x"20616363",
001454 => x"6573733A",
001455 => x"20000000",
001456 => x"210A0D00",
001457 => x"446F6E65",
001458 => x"204C6F61",
001459 => x"64696E67",
001460 => x"210D0A00",
001461 => x"4C415354",
001462 => x"20414444",
001463 => x"52455353",
001464 => x"3A000000",
001465 => x"20496E76",
001466 => x"616C6964",
001467 => x"2070726F",
001468 => x"6772616D",
001469 => x"6D696E67",
001470 => x"2066696C",
001471 => x"65210D0A",
001472 => x"0D0A5365",
001473 => x"6C656374",
001474 => x"3A200000",
001475 => x"0D0A0D0A",
001476 => x"41626F72",
001477 => x"74206475",
001478 => x"6D70696E",
001479 => x"67206279",
001480 => x"20707265",
001481 => x"7373696E",
001482 => x"6720616E",
001483 => x"79206B65",
001484 => x"792E0D0A",
001485 => x"50726573",
001486 => x"7320616E",
001487 => x"79206B65",
001488 => x"7920746F",
001489 => x"20636F6E",
001490 => x"74696E75",
001491 => x"652E0D0A",
001492 => x"0D0A0000",
001493 => x"0D0A0D0A",
001494 => x"44756D70",
001495 => x"696E6720",
001496 => x"636F6D70",
001497 => x"6C657465",
001498 => x"642E0D0A",
001499 => x"0D0A5365",
001500 => x"6C656374",
001501 => x"3A200000",
001502 => x"0D0A0D0A",
001503 => x"456E7465",
001504 => x"72206465",
001505 => x"76696365",
001506 => x"20616464",
001507 => x"72657373",
001508 => x"20283278",
001509 => x"20686578",
001510 => x"5F636861",
001511 => x"72732C20",
001512 => x"73657420",
001513 => x"4C534220",
001514 => x"746F2027",
001515 => x"3027293A",
001516 => x"20000000",
001517 => x"20496E76",
001518 => x"616C6964",
001519 => x"20616464",
001520 => x"72657373",
001521 => x"210D0A0D",
001522 => x"0A53656C",
001523 => x"6563743A",
001524 => x"20000000",
001525 => x"0D0A4170",
001526 => x"706C6963",
001527 => x"6174696F",
001528 => x"6E207769",
001529 => x"6C6C2073",
001530 => x"74617274",
001531 => x"20617574",
001532 => x"6F6D6174",
001533 => x"6963616C",
001534 => x"6C792061",
001535 => x"66746572",
001536 => x"2075706C",
001537 => x"6F61642E",
001538 => x"0D0A2D3E",
001539 => x"204C6F61",
001540 => x"64696E67",
001541 => x"20626F6F",
001542 => x"7420696D",
001543 => x"6167652E",
001544 => x"2E2E0000",
001545 => x"2055706C",
001546 => x"6F616420",
001547 => x"636F6D70",
001548 => x"6C657465",
001549 => x"0D0A0000",
001550 => x"20496E76",
001551 => x"616C6964",
001552 => x"20626F6F",
001553 => x"74206465",
001554 => x"76696365",
001555 => x"206F7220",
001556 => x"66696C65",
001557 => x"210D0A0D",
001558 => x"0A53656C",
001559 => x"6563743A",
001560 => x"20000000",
001561 => x"0D0A496E",
001562 => x"76616C69",
001563 => x"64206164",
001564 => x"64726573",
001565 => x"73210D0A",
001566 => x"0D0A5365",
001567 => x"6C656374",
001568 => x"3A200000",
001569 => x"0D0A4461",
001570 => x"74612077",
001571 => x"696C6C20",
001572 => x"6F766572",
001573 => x"77726974",
001574 => x"65205241",
001575 => x"4D20636F",
001576 => x"6E74656E",
001577 => x"74210D0A",
001578 => x"2D3E2057",
001579 => x"61697469",
001580 => x"6E672066",
001581 => x"6F722027",
001582 => x"73746F72",
001583 => x"6D5F7072",
001584 => x"6F677261",
001585 => x"6D2E6269",
001586 => x"6E272069",
001587 => x"6E206279",
001588 => x"74652D73",
001589 => x"74726561",
001590 => x"6D206D6F",
001591 => x"64652E2E",
001592 => x"2E000000",
001593 => x"20455252",
001594 => x"4F522120",
001595 => x"50726F67",
001596 => x"72616D20",
001597 => x"66696C65",
001598 => x"20746F6F",
001599 => x"20626967",
001600 => x"210D0A0D",
001601 => x"0A000000",
001602 => x"20446F77",
001603 => x"6E6C6F61",
001604 => x"6420636F",
001605 => x"6D706C65",
001606 => x"7465640D",
001607 => x"0A000000",
001608 => x"57726974",
001609 => x"696E6720",
001610 => x"62756666",
001611 => x"65722074",
001612 => x"6F206932",
001613 => x"63204545",
001614 => x"50524F4D",
001615 => x"2E2E2E00",
001616 => x"20436F6D",
001617 => x"706C6574",
001618 => x"65640D0A",
001619 => x"0D0A0000",
001620 => x"20496E76",
001621 => x"616C6964",
001622 => x"20626F6F",
001623 => x"74206465",
001624 => x"76696365",
001625 => x"206F7220",
001626 => x"66696C65",
001627 => x"210D0A0D",
001628 => x"0A000000",
001629 => x"0D0A0D0A",
001630 => x"456E7465",
001631 => x"72206465",
001632 => x"76696365",
001633 => x"20616464",
001634 => x"72657373",
001635 => x"20283220",
001636 => x"6865782D",
001637 => x"63686172",
001638 => x"732C2073",
001639 => x"6574204C",
001640 => x"53422074",
001641 => x"6F202730",
001642 => x"27293A20",
001643 => x"00000000",
001644 => x"0D0A0D0A",
001645 => x"41626F72",
001646 => x"74206475",
001647 => x"6D70696E",
001648 => x"67206279",
001649 => x"20707265",
001650 => x"7373696E",
001651 => x"6720616E",
001652 => x"79206B65",
001653 => x"792E2049",
001654 => x"66206E6F",
001655 => x"20646174",
001656 => x"61206973",
001657 => x"2073686F",
001658 => x"776E2C0D",
001659 => x"0A000000",
001660 => x"74686520",
001661 => x"73656C65",
001662 => x"63746564",
001663 => x"20646576",
001664 => x"69636520",
001665 => x"6973206E",
001666 => x"6F742072",
001667 => x"6573706F",
001668 => x"6E64696E",
001669 => x"672E2050",
001670 => x"72657373",
001671 => x"20616E79",
001672 => x"206B6579",
001673 => x"20746F20",
001674 => x"636F6E74",
001675 => x"696E7565",
001676 => x"2E0D0A0D",
001677 => x"0A000000",
001678 => x"0D0A0D0A",
001679 => x"4175746F",
001680 => x"6D617469",
001681 => x"6320626F",
001682 => x"6F742063",
001683 => x"6F6E6669",
001684 => x"67757261",
001685 => x"74696F6E",
001686 => x"20666F72",
001687 => x"20706F77",
001688 => x"65722D75",
001689 => x"703A0D0A",
001690 => x"00000000",
001691 => x"5B333231",
001692 => x"305D2063",
001693 => x"6F6E6669",
001694 => x"67757261",
001695 => x"74696F6E",
001696 => x"20444950",
001697 => x"20737769",
001698 => x"7463680D",
001699 => x"0A203030",
001700 => x"3030202D",
001701 => x"20537461",
001702 => x"72742062",
001703 => x"6F6F746C",
001704 => x"6F616465",
001705 => x"7220636F",
001706 => x"6E736F6C",
001707 => x"650D0A20",
001708 => x"30303031",
001709 => x"202D2041",
001710 => x"75746F6D",
001711 => x"61746963",
001712 => x"20626F6F",
001713 => x"74206672",
001714 => x"6F6D2063",
001715 => x"6F726520",
001716 => x"52414D0D",
001717 => x"0A000000",
001718 => x"20303031",
001719 => x"30202D20",
001720 => x"4175746F",
001721 => x"6D617469",
001722 => x"6320626F",
001723 => x"6F742066",
001724 => x"726F6D20",
001725 => x"49324320",
001726 => x"45455052",
001727 => x"4F4D2028",
001728 => x"41646472",
001729 => x"65737320",
001730 => x"30784130",
001731 => x"290D0A0D",
001732 => x"0A53656C",
001733 => x"6563743A",
001734 => x"20000000",
001735 => x"0D0A0D0A",
001736 => x"5765276C",
001737 => x"6C207365",
001738 => x"6E642079",
001739 => x"6F752062",
001740 => x"61636B20",
001741 => x"2D20746F",
001742 => x"20746865",
001743 => x"20667574",
001744 => x"75726521",
001745 => x"2E0D0A0D",
001746 => x"0A000000",
001747 => x"202D2044",
001748 => x"6F63746F",
001749 => x"7220456D",
001750 => x"6D657420",
001751 => x"4C2E2042",
001752 => x"726F776E",
001753 => x"0D0A0D0A",
001754 => x"53656C65",
001755 => x"63743A20",
001756 => x"00000000",
001757 => x"20496E76",
001758 => x"616C6964",
001759 => x"206F7065",
001760 => x"72617469",
001761 => x"6F6E210D",
001762 => x"0A547279",
001763 => x"20616761",
001764 => x"696E3A20",
001765 => x"00000000",
001766 => x"0D0A0D0A",
001767 => x"2D3E2053",
001768 => x"74617274",
001769 => x"696E6720",
001770 => x"6170706C",
001771 => x"69636174",
001772 => x"696F6E2E",
001773 => x"2E2E0D0A",
001774 => x"0D0A0000",
001775 => x"0D0A0D0A",
001776 => x"2D3E2064",
001777 => x"69736162",
001778 => x"6C652077",
001779 => x"72697465",
001780 => x"2D746872",
001781 => x"6F756768",
001782 => x"20737472",
001783 => x"61746567",
001784 => x"792E2E2E",
001785 => x"0D0A0D0A",
001786 => x"00000000",
001787 => x"0D0A0D0A",
001788 => x"2D3E206A",
001789 => x"756D7020",
001790 => x"746F2061",
001791 => x"70706C69",
001792 => x"63617469",
001793 => x"6F6E2E2E",
001794 => x"2E0D0A0D",
001795 => x"0A000000",
001796 => x"21217368",
001797 => x"6F756C64",
001798 => x"206E6F74",
001799 => x"20626520",
001800 => x"68657265",
001801 => x"21210D0A",
001802 => x"00000000",
001803 => x"0D0A0D0A",
001804 => x"41626F72",
001805 => x"74656421",
001806 => x"00000000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;