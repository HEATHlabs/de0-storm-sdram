-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
	--regular bootloader
000000 => x"EA000006",
000001 => x"EAFFFFFE",
000002 => x"EAFFFFFE",
000003 => x"EAFFFFFE",
000004 => x"EAFFFFFE",
000005 => x"E1A00000",
000006 => x"EAFFFFFE",
000007 => x"EAFFFFFE",
000008 => x"E59F0040",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA018",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"E1A04000",
000023 => x"E3A00000",
000024 => x"E1A0F004",
000025 => x"EAFFFFFE",
000026 => x"00002000",
000027 => x"000107BC",
000028 => x"E3E03A0F",
000029 => x"E5131FFB",
000030 => x"E20020FF",
000031 => x"E3A00001",
000032 => x"E0010210",
000033 => x"E1A0F00E",
000034 => x"E3E03A0F",
000035 => x"E5130FFB",
000036 => x"E1A0F00E",
000037 => x"E3E01A0F",
000038 => x"E5113FFF",
000039 => x"E20000FF",
000040 => x"E3A02001",
000041 => x"E1833012",
000042 => x"E5013FFF",
000043 => x"E1A0F00E",
000044 => x"E20000FF",
000045 => x"E3A02001",
000046 => x"E1A02012",
000047 => x"E3E01A0F",
000048 => x"E5113FFF",
000049 => x"E1E02002",
000050 => x"E0033002",
000051 => x"E5013FFF",
000052 => x"E1A0F00E",
000053 => x"E3E01A0F",
000054 => x"E5113FFF",
000055 => x"E20000FF",
000056 => x"E3A02001",
000057 => x"E0233012",
000058 => x"E5013FFF",
000059 => x"E1A0F00E",
000060 => x"E3E03A0F",
000061 => x"E5030FFF",
000062 => x"E1A0F00E",
000063 => x"E20000FF",
000064 => x"E3500007",
000065 => x"E92D4010",
000066 => x"E3A0C000",
000067 => x"E3E0E0FF",
000068 => x"E20110FF",
000069 => x"8A000011",
000070 => x"E2403004",
000071 => x"E20330FF",
000072 => x"E3500003",
000073 => x"E1A0E183",
000074 => x"E3E04A0F",
000075 => x"E1A0C180",
000076 => x"9A000007",
000077 => x"E3A030FF",
000078 => x"E1A03E13",
000079 => x"E5142F8B",
000080 => x"E1E03003",
000081 => x"E0022003",
000082 => x"E1822E11",
000083 => x"E5042F8B",
000084 => x"E8BD8010",
000085 => x"E3A030FF",
000086 => x"E1A03C13",
000087 => x"E1E0E003",
000088 => x"E3E02A0F",
000089 => x"E5123F8F",
000090 => x"E003300E",
000091 => x"E1833C11",
000092 => x"E5023F8F",
000093 => x"E8BD8010",
000094 => x"E20000FF",
000095 => x"E3500007",
000096 => x"E3A02000",
000097 => x"8A00000A",
000098 => x"E2403004",
000099 => x"E3500003",
000100 => x"E20320FF",
000101 => x"9A000005",
000102 => x"E3E03A0F",
000103 => x"E5130F8B",
000104 => x"E1A02182",
000105 => x"E1A00230",
000106 => x"E20000FF",
000107 => x"E1A0F00E",
000108 => x"E1A02180",
000109 => x"E3E03A0F",
000110 => x"E5130F8F",
000111 => x"E1A00230",
000112 => x"E20000FF",
000113 => x"E1A0F00E",
000114 => x"E3E02A0F",
000115 => x"E5123EFB",
000116 => x"E3130002",
000117 => x"E3E00000",
000118 => x"15120EFF",
000119 => x"E1A0F00E",
000120 => x"E3E02A0F",
000121 => x"E5123EFB",
000122 => x"E3130001",
000123 => x"0AFFFFFC",
000124 => x"E20030FF",
000125 => x"E5023EFF",
000126 => x"E1A0F00E",
000127 => x"E20000FF",
000128 => x"E3500001",
000129 => x"E3812B01",
000130 => x"03E03A0F",
000131 => x"E3811B09",
000132 => x"13E03A0F",
000133 => x"05031CFF",
000134 => x"15032CFF",
000135 => x"E1A0F00E",
000136 => x"E3E03A0F",
000137 => x"E5030CFB",
000138 => x"E1A0F00E",
000139 => x"E3E02A0F",
000140 => x"E5123CFF",
000141 => x"E3130C01",
000142 => x"1AFFFFFC",
000143 => x"E5020CEF",
000144 => x"E5123CFF",
000145 => x"E3833C01",
000146 => x"E5023CFF",
000147 => x"E3E02A0F",
000148 => x"E5123CFF",
000149 => x"E3130C01",
000150 => x"1AFFFFFC",
000151 => x"E5120CEF",
000152 => x"E1A0F00E",
000153 => x"E3E01A0F",
000154 => x"E5113CF7",
000155 => x"E20000FF",
000156 => x"E3A02001",
000157 => x"E1833012",
000158 => x"E5013CF7",
000159 => x"E1A0F00E",
000160 => x"E20000FF",
000161 => x"E3A02001",
000162 => x"E1A02012",
000163 => x"E3E01A0F",
000164 => x"E5113CF7",
000165 => x"E1E02002",
000166 => x"E0033002",
000167 => x"E5013CF7",
000168 => x"E1A0F00E",
000169 => x"E3E02A0F",
000170 => x"E5123BE7",
000171 => x"E1A01420",
000172 => x"E3C33080",
000173 => x"E5023BE7",
000174 => x"E5020BEF",
000175 => x"E5021BEB",
000176 => x"E5123BE7",
000177 => x"E3833080",
000178 => x"E5023BE7",
000179 => x"E1A0F00E",
000180 => x"E92D4030",
000181 => x"E3A0C090",
000182 => x"E20140FE",
000183 => x"E3E0EA0F",
000184 => x"E5DD500F",
000185 => x"E20000FF",
000186 => x"E50E4BE3",
000187 => x"E20110FF",
000188 => x"E50ECBFF",
000189 => x"E1A04002",
000190 => x"E203C0FF",
000191 => x"E51E3BFF",
000192 => x"E3130002",
000193 => x"1AFFFFFC",
000194 => x"E51E3BFF",
000195 => x"E3130080",
000196 => x"13E00000",
000197 => x"18BD8030",
000198 => x"E35C0000",
000199 => x"0A000012",
000200 => x"E24C3001",
000201 => x"E203C0FF",
000202 => x"E35C0001",
000203 => x"01A02424",
000204 => x"03E03A0F",
000205 => x"13E03A0F",
000206 => x"05032BE3",
000207 => x"15034BE3",
000208 => x"E3E02A0F",
000209 => x"E3A03010",
000210 => x"E5023BFF",
000211 => x"E5123BFF",
000212 => x"E3130002",
000213 => x"1AFFFFFC",
000214 => x"E5123BFF",
000215 => x"E3130080",
000216 => x"0AFFFFEC",
000217 => x"E3E00001",
000218 => x"E8BD8030",
000219 => x"E3500077",
000220 => x"1A00000C",
000221 => x"E3E03A0F",
000222 => x"E3A02050",
000223 => x"E5035BE3",
000224 => x"E5032BFF",
000225 => x"E1A02003",
000226 => x"E5123BFF",
000227 => x"E3130002",
000228 => x"1AFFFFFC",
000229 => x"E5123BFF",
000230 => x"E2130080",
000231 => x"08BD8030",
000232 => x"E3E00002",
000233 => x"E8BD8030",
000234 => x"E3500072",
000235 => x"13E00003",
000236 => x"18BD8030",
000237 => x"E3813001",
000238 => x"E3E02A0F",
000239 => x"E3A01090",
000240 => x"E5023BE3",
000241 => x"E5021BFF",
000242 => x"E5123BFF",
000243 => x"E3130002",
000244 => x"1AFFFFFC",
000245 => x"E5123BFF",
000246 => x"E3130080",
000247 => x"1AFFFFEF",
000248 => x"E3A03068",
000249 => x"E5023BFF",
000250 => x"E3E00A0F",
000251 => x"E5103BFF",
000252 => x"E3130002",
000253 => x"1AFFFFFC",
000254 => x"E5100BE3",
000255 => x"E8BD8030",
000256 => x"E20000FF",
000257 => x"E350000F",
000258 => x"979FF100",
000259 => x"EA00000F",
000260 => x"000104D0",
000261 => x"000104C8",
000262 => x"000104C0",
000263 => x"000104B8",
000264 => x"000104B0",
000265 => x"000104A8",
000266 => x"000104A0",
000267 => x"00010498",
000268 => x"00010490",
000269 => x"00010488",
000270 => x"00010480",
000271 => x"00010478",
000272 => x"00010470",
000273 => x"00010468",
000274 => x"00010460",
000275 => x"00010458",
000276 => x"E3A00000",
000277 => x"E1A0F00E",
000278 => x"EE1F0F1F",
000279 => x"E1A0F00E",
000280 => x"EE1E0F1E",
000281 => x"E1A0F00E",
000282 => x"EE1D0F1D",
000283 => x"E1A0F00E",
000284 => x"EE1C0F1C",
000285 => x"E1A0F00E",
000286 => x"EE1B0F1B",
000287 => x"E1A0F00E",
000288 => x"EE1A0F1A",
000289 => x"E1A0F00E",
000290 => x"EE190F19",
000291 => x"E1A0F00E",
000292 => x"EE180F18",
000293 => x"E1A0F00E",
000294 => x"EE170F17",
000295 => x"E1A0F00E",
000296 => x"EE160F16",
000297 => x"E1A0F00E",
000298 => x"EE150F15",
000299 => x"E1A0F00E",
000300 => x"EE140F14",
000301 => x"E1A0F00E",
000302 => x"EE130F13",
000303 => x"E1A0F00E",
000304 => x"EE120F12",
000305 => x"E1A0F00E",
000306 => x"EE110F11",
000307 => x"E1A0F00E",
000308 => x"EE100F10",
000309 => x"E1A0F00E",
000310 => x"E20110FF",
000311 => x"E2411006",
000312 => x"E3510007",
000313 => x"979FF101",
000314 => x"EA000008",
000315 => x"00010514",
000316 => x"00010510",
000317 => x"00010510",
000318 => x"00010510",
000319 => x"00010510",
000320 => x"0001051C",
000321 => x"00010524",
000322 => x"0001050C",
000323 => x"EE0D0F1D",
000324 => x"E1A0F00E",
000325 => x"EE060F16",
000326 => x"E1A0F00E",
000327 => x"EE0B0F1B",
000328 => x"E1A0F00E",
000329 => x"EE0C0F1C",
000330 => x"E1A0F00E",
000331 => x"E92D4010",
000332 => x"E1A04000",
000333 => x"E5D00000",
000334 => x"E3500000",
000335 => x"1A000003",
000336 => x"EA000005",
000337 => x"E5F40001",
000338 => x"E3500000",
000339 => x"0A000002",
000340 => x"EBFFFF22",
000341 => x"E3500000",
000342 => x"CAFFFFF9",
000343 => x"E1A00004",
000344 => x"E8BD8010",
000345 => x"E92D4070",
000346 => x"E2514000",
000347 => x"E1A05000",
000348 => x"E20260FF",
000349 => x"DA00000B",
000350 => x"EBFFFF12",
000351 => x"E3700001",
000352 => x"E20030FF",
000353 => x"0A000005",
000354 => x"E3560001",
000355 => x"E5C53000",
000356 => x"E1A00003",
000357 => x"E2855001",
000358 => x"0A000005",
000359 => x"E2444001",
000360 => x"E3540000",
000361 => x"CAFFFFF3",
000362 => x"E59F300C",
000363 => x"E5C53000",
000364 => x"E8BD8070",
000365 => x"EBFFFF09",
000366 => x"EAFFFFF7",
000367 => x"000111A4",
000368 => x"E92D4030",
000369 => x"E2514000",
000370 => x"E1A05000",
000371 => x"D8BD8030",
000372 => x"E4D50001",
000373 => x"EBFFFF01",
000374 => x"E2544001",
000375 => x"1AFFFFFB",
000376 => x"E8BD8030",
000377 => x"E92D4010",
000378 => x"E20240FF",
000379 => x"E3540008",
000380 => x"83A04008",
000381 => x"8A000001",
000382 => x"E3540000",
000383 => x"03A04001",
000384 => x"E1A02001",
000385 => x"E1A0E004",
000386 => x"E1A0310E",
000387 => x"E35E0001",
000388 => x"E2433004",
000389 => x"E1A0C000",
000390 => x"81A0C330",
000391 => x"E24E3001",
000392 => x"E20CC00F",
000393 => x"E203E0FF",
000394 => x"E35C0009",
000395 => x"E28C3030",
000396 => x"828C3037",
000397 => x"E35E0000",
000398 => x"E4C23001",
000399 => x"1AFFFFF1",
000400 => x"E2443001",
000401 => x"E20330FF",
000402 => x"E0813003",
000403 => x"E5C3E001",
000404 => x"E8BD8010",
000405 => x"E92D4010",
000406 => x"E1A04000",
000407 => x"E3540007",
000408 => x"E3A01010",
000409 => x"E3A00001",
000410 => x"9A000001",
000411 => x"E3A00000",
000412 => x"E8BD8010",
000413 => x"EBFFFEE0",
000414 => x"E3A00006",
000415 => x"EBFFFEF8",
000416 => x"E3A00000",
000417 => x"EBFFFEE8",
000418 => x"E1A00584",
000419 => x"E8BD4010",
000420 => x"EAFFFEE5",
000421 => x"E0603280",
000422 => x"E0800103",
000423 => x"E0800100",
000424 => x"E1A00200",
000425 => x"E3500000",
000426 => x"D1A0F00E",
000427 => x"E1A00000",
000428 => x"E2500001",
000429 => x"1AFFFFFC",
000430 => x"E1A0F00E",
000431 => x"E212C0FF",
000432 => x"0A00000B",
000433 => x"E5D02000",
000434 => x"E5D13000",
000435 => x"E1520003",
000436 => x"0A000004",
000437 => x"EA000008",
000438 => x"E5F02001",
000439 => x"E5F13001",
000440 => x"E1520003",
000441 => x"1A000004",
000442 => x"E24C3001",
000443 => x"E213C0FF",
000444 => x"1AFFFFF8",
000445 => x"E3A00001",
000446 => x"E1A0F00E",
000447 => x"E3A00000",
000448 => x"E1A0F00E",
000449 => x"E92D4030",
000450 => x"E1A04081",
000451 => x"E3540000",
000452 => x"E1A05000",
000453 => x"D3A00000",
000454 => x"D8BD8030",
000455 => x"E3A00000",
000456 => x"E1A01000",
000457 => x"E7D12005",
000458 => x"E2423030",
000459 => x"E082C200",
000460 => x"E3530009",
000461 => x"E242E041",
000462 => x"924C0030",
000463 => x"9A000007",
000464 => x"E0823200",
000465 => x"E35E0005",
000466 => x"E242C061",
000467 => x"92430037",
000468 => x"9A000002",
000469 => x"E0823200",
000470 => x"E35C0005",
000471 => x"92430057",
000472 => x"E2811001",
000473 => x"E1510004",
000474 => x"1AFFFFED",
000475 => x"E8BD8030",
000476 => x"E5D03003",
000477 => x"E5D02002",
000478 => x"E5D01000",
000479 => x"E1833402",
000480 => x"E5D00001",
000481 => x"E1833C01",
000482 => x"E1830800",
000483 => x"E1A0F00E",
000484 => x"E52DE004",
000485 => x"E59F0014",
000486 => x"EBFFFF63",
000487 => x"E59F0010",
000488 => x"EBFFFF61",
000489 => x"E59F000C",
000490 => x"E49DE004",
000491 => x"EAFFFF5E",
000492 => x"000111A8",
000493 => x"0001120C",
000494 => x"00011270",
000495 => x"E92D45F0",
000496 => x"E3A00000",
000497 => x"E24DD014",
000498 => x"EBFFFE48",
000499 => x"E3A0100D",
000500 => x"E3A000C3",
000501 => x"EBFFFF3F",
000502 => x"E3A00063",
000503 => x"EBFFFEB0",
000504 => x"E3A00006",
000505 => x"EBFFFF05",
000506 => x"E3A01006",
000507 => x"E3800008",
000508 => x"EBFFFF38",
000509 => x"E3A0000D",
000510 => x"EBFFFF00",
000511 => x"E1A008A0",
000512 => x"E1E00000",
000513 => x"E200000F",
000514 => x"E3500001",
000515 => x"03A04030",
000516 => x"028DA00F",
000517 => x"0A000020",
000518 => x"E3500002",
000519 => x"0A00008C",
000520 => x"E59F0874",
000521 => x"EBFFFF40",
000522 => x"E59F0870",
000523 => x"EBFFFF3E",
000524 => x"E59F086C",
000525 => x"EBFFFF3C",
000526 => x"E59F0868",
000527 => x"EBFFFF3A",
000528 => x"E59F0864",
000529 => x"EBFFFF38",
000530 => x"E59F0860",
000531 => x"EBFFFF36",
000532 => x"E59F085C",
000533 => x"EBFFFF34",
000534 => x"E59F0858",
000535 => x"EBFFFF32",
000536 => x"E28D4006",
000537 => x"E59F0850",
000538 => x"EBFFFF2F",
000539 => x"E1A01004",
000540 => x"E3A02008",
000541 => x"E3A00401",
000542 => x"EBFFFF59",
000543 => x"E1A00004",
000544 => x"EBFFFF29",
000545 => x"E59F0834",
000546 => x"EBFFFF27",
000547 => x"EBFFFFBF",
000548 => x"E28DA00F",
000549 => x"EBFFFE4B",
000550 => x"E1A04000",
000551 => x"E3A0000D",
000552 => x"EBFFFED6",
000553 => x"E3100801",
000554 => x"03A06001",
000555 => x"03A050A0",
000556 => x"1A00004B",
000557 => x"E3A04000",
000558 => x"E59F0804",
000559 => x"EBFFFF1A",
000560 => x"E1A01005",
000561 => x"E1A02004",
000562 => x"E3A03002",
000563 => x"E3A00072",
000564 => x"E58D4000",
000565 => x"EBFFFE7D",
000566 => x"E1A01005",
000567 => x"E5CD000F",
000568 => x"E3A02001",
000569 => x"E3A03002",
000570 => x"E3A00072",
000571 => x"E58D4000",
000572 => x"EBFFFE76",
000573 => x"E3A02002",
000574 => x"E1A03002",
000575 => x"E5CD0010",
000576 => x"E1A01005",
000577 => x"E3A00072",
000578 => x"E58D4000",
000579 => x"EBFFFE6F",
000580 => x"E3A03002",
000581 => x"E5CD0011",
000582 => x"E1A01005",
000583 => x"E3A00072",
000584 => x"E3A02003",
000585 => x"E58D4000",
000586 => x"EBFFFE68",
000587 => x"E5DD300F",
000588 => x"E20000FF",
000589 => x"E3530053",
000590 => x"E5CD0012",
000591 => x"1A000002",
000592 => x"E5DD3010",
000593 => x"E353004D",
000594 => x"0A000078",
000595 => x"E59F0774",
000596 => x"EBFFFEF5",
000597 => x"E3560000",
000598 => x"0AFFFFCD",
000599 => x"E59F0768",
000600 => x"EBFFFEF1",
000601 => x"E3A0100D",
000602 => x"E3A00000",
000603 => x"EBFFFED9",
000604 => x"E3A00006",
000605 => x"EBFFFEA1",
000606 => x"E3A01006",
000607 => x"E3C00008",
000608 => x"EBFFFED4",
000609 => x"E3A00006",
000610 => x"EBFFFE9C",
000611 => x"E1E00000",
000612 => x"E2000002",
000613 => x"E3A01006",
000614 => x"E1E00000",
000615 => x"EBFFFECD",
000616 => x"E3A00006",
000617 => x"EBFFFE95",
000618 => x"E1E00000",
000619 => x"E2000004",
000620 => x"E3A01006",
000621 => x"E1E00000",
000622 => x"EBFFFEC6",
000623 => x"E3A00006",
000624 => x"EBFFFE8E",
000625 => x"E1A00800",
000626 => x"E1A00820",
000627 => x"E3800702",
000628 => x"E3A01006",
000629 => x"EBFFFEBF",
000630 => x"E3A00401",
000631 => x"EBFFFD9D",
000632 => x"EAFFFFFE",
000633 => x"E3540034",
000634 => x"0A000028",
000635 => x"CA00001B",
000636 => x"E3540031",
000637 => x"0A000035",
000638 => x"DA000097",
000639 => x"E3540032",
000640 => x"0A0000A1",
000641 => x"E3540033",
000642 => x"1A000097",
000643 => x"E1A00004",
000644 => x"EBFFFDF2",
000645 => x"E59F06B4",
000646 => x"EBFFFEC3",
000647 => x"E1A0000A",
000648 => x"E3A01002",
000649 => x"E3A02001",
000650 => x"EBFFFECD",
000651 => x"E3A01002",
000652 => x"E1A0000A",
000653 => x"EBFFFF32",
000654 => x"E21010FF",
000655 => x"11A05001",
000656 => x"13A06000",
000657 => x"1AFFFF9A",
000658 => x"E59F0684",
000659 => x"EBFFFEB6",
000660 => x"EAFFFF8F",
000661 => x"E3A04033",
000662 => x"E28DA00F",
000663 => x"EAFFFF8E",
000664 => x"E3540066",
000665 => x"0A00002A",
000666 => x"DA0000A8",
000667 => x"E3540068",
000668 => x"0A00010A",
000669 => x"E3540072",
000670 => x"1A00007B",
000671 => x"E1A00004",
000672 => x"EBFFFDD6",
000673 => x"E3A006FF",
000674 => x"E280F20F",
000675 => x"EAFFFFFE",
000676 => x"E1A00004",
000677 => x"EBFFFDD1",
000678 => x"E59F0630",
000679 => x"EBFFFEA2",
000680 => x"E1A0000A",
000681 => x"E3A01002",
000682 => x"E3A02001",
000683 => x"EBFFFEAC",
000684 => x"E1A0000A",
000685 => x"E3A01002",
000686 => x"EBFFFF11",
000687 => x"E21080FF",
000688 => x"1A00009F",
000689 => x"E59F060C",
000690 => x"EBFFFE97",
000691 => x"EAFFFF70",
000692 => x"E1A00004",
000693 => x"EBFFFDC1",
000694 => x"E59F05FC",
000695 => x"EBFFFE92",
000696 => x"E1A0000A",
000697 => x"E3A01004",
000698 => x"E3A02000",
000699 => x"EBFFFE9C",
000700 => x"E5DD300F",
000701 => x"E3530053",
000702 => x"1A000002",
000703 => x"E5DD3010",
000704 => x"E353004D",
000705 => x"0A000110",
000706 => x"E59F05D0",
000707 => x"EBFFFE86",
000708 => x"EAFFFF5F",
000709 => x"E1A00004",
000710 => x"EBFFFDB0",
000711 => x"E59F05C0",
000712 => x"EBFFFE81",
000713 => x"E59F05BC",
000714 => x"EBFFFE7F",
000715 => x"EAFFFF58",
000716 => x"E5DD3011",
000717 => x"E3530042",
000718 => x"1AFFFF83",
000719 => x"E3500052",
000720 => x"1AFFFF81",
000721 => x"E1A01005",
000722 => x"E3A02004",
000723 => x"E2433040",
000724 => x"E2800020",
000725 => x"E58D4000",
000726 => x"EBFFFDDC",
000727 => x"E1A01005",
000728 => x"E5CD000F",
000729 => x"E3A02005",
000730 => x"E3A03002",
000731 => x"E3A00072",
000732 => x"E58D4000",
000733 => x"EBFFFDD5",
000734 => x"E1A01005",
000735 => x"E5CD0010",
000736 => x"E3A02006",
000737 => x"E3A03002",
000738 => x"E3A00072",
000739 => x"E58D4000",
000740 => x"EBFFFDCE",
000741 => x"E1A01005",
000742 => x"E5CD0011",
000743 => x"E3A02007",
000744 => x"E3A03002",
000745 => x"E3A00072",
000746 => x"E58D4000",
000747 => x"EBFFFDC7",
000748 => x"E5CD0012",
000749 => x"E1A0000A",
000750 => x"EBFFFEEC",
000751 => x"E2907004",
000752 => x"0A000022",
000753 => x"E1A06004",
000754 => x"E2842008",
000755 => x"E1A01005",
000756 => x"E3A03002",
000757 => x"E3A00072",
000758 => x"E58D6000",
000759 => x"EBFFFDBB",
000760 => x"E2842009",
000761 => x"E5CD000F",
000762 => x"E1A01005",
000763 => x"E3A03002",
000764 => x"E3A00072",
000765 => x"E58D6000",
000766 => x"EBFFFDB4",
000767 => x"E284200A",
000768 => x"E5CD0010",
000769 => x"E1A01005",
000770 => x"E3A03002",
000771 => x"E3A00072",
000772 => x"E58D6000",
000773 => x"EBFFFDAD",
000774 => x"E284200B",
000775 => x"E5CD0011",
000776 => x"E1A01005",
000777 => x"E3A03002",
000778 => x"E3A00072",
000779 => x"E58D6000",
000780 => x"EBFFFDA6",
000781 => x"E5CD0012",
000782 => x"E1A0000A",
000783 => x"EBFFFECB",
000784 => x"E4840004",
000785 => x"E1540007",
000786 => x"13540902",
000787 => x"3AFFFFDD",
000788 => x"E59F0494",
000789 => x"EBFFFE34",
000790 => x"EAFFFF3F",
000791 => x"E3740001",
000792 => x"0AFFFF0B",
000793 => x"E3540030",
000794 => x"0A000004",
000795 => x"E20400FF",
000796 => x"EBFFFD5A",
000797 => x"E59F0474",
000798 => x"EBFFFE2B",
000799 => x"EAFFFF04",
000800 => x"E1A00004",
000801 => x"EBFFFD55",
000802 => x"EAFFFF33",
000803 => x"E1A00004",
000804 => x"EBFFFD52",
000805 => x"E59F0458",
000806 => x"EBFFFE23",
000807 => x"EBFFFD49",
000808 => x"E3700001",
000809 => x"0AFFFFFC",
000810 => x"EBFFFD46",
000811 => x"E3700001",
000812 => x"1AFFFFFC",
000813 => x"E3A05401",
000814 => x"EA000001",
000815 => x"E1550003",
000816 => x"0A00000F",
000817 => x"E5954000",
000818 => x"E1A00C24",
000819 => x"EBFFFD43",
000820 => x"E1A00824",
000821 => x"EBFFFD41",
000822 => x"E1A00424",
000823 => x"EBFFFD3F",
000824 => x"E1A00004",
000825 => x"EBFFFD3D",
000826 => x"EBFFFD36",
000827 => x"E3A03401",
000828 => x"E2833E9E",
000829 => x"E3700001",
000830 => x"E2855004",
000831 => x"E2833004",
000832 => x"0AFFFFED",
000833 => x"E59F03EC",
000834 => x"EBFFFE07",
000835 => x"EAFFFEE0",
000836 => x"E3540035",
000837 => x"0A0000AC",
000838 => x"E3540061",
000839 => x"1AFFFFD2",
000840 => x"E1A00004",
000841 => x"EBFFFD2D",
000842 => x"E59F03CC",
000843 => x"EBFFFDFE",
000844 => x"E59F03C8",
000845 => x"EBFFFDFC",
000846 => x"E59F03C4",
000847 => x"EBFFFDFA",
000848 => x"EAFFFED3",
000849 => x"E59F03BC",
000850 => x"EBFFFDF7",
000851 => x"E1A0000A",
000852 => x"E3A01004",
000853 => x"E3A02000",
000854 => x"EBFFFE01",
000855 => x"E5DD300F",
000856 => x"E3530053",
000857 => x"1A000002",
000858 => x"E5DD2010",
000859 => x"E352004D",
000860 => x"0A000004",
000861 => x"E59F0390",
000862 => x"EBFFFDEB",
000863 => x"E59F038C",
000864 => x"EBFFFDE9",
000865 => x"EAFFFEC2",
000866 => x"E5DD1011",
000867 => x"E3510042",
000868 => x"1AFFFFF7",
000869 => x"E5DD0012",
000870 => x"E3500052",
000871 => x"1AFFFFF4",
000872 => x"E3A04000",
000873 => x"E5C43000",
000874 => x"E1A00000",
000875 => x"E5C42001",
000876 => x"E1A00000",
000877 => x"E5C41002",
000878 => x"E1A00000",
000879 => x"E5C40003",
000880 => x"E1A00000",
000881 => x"E241103E",
000882 => x"E1A0000A",
000883 => x"E1A02004",
000884 => x"EBFFFDE3",
000885 => x"E5DD300F",
000886 => x"E5C43004",
000887 => x"E5DD2010",
000888 => x"E5C42005",
000889 => x"E5DD3011",
000890 => x"E5C43006",
000891 => x"E5DD2012",
000892 => x"E1A0000A",
000893 => x"E5C42007",
000894 => x"EBFFFE5C",
000895 => x"E3A03CFF",
000896 => x"E28330FC",
000897 => x"E1500003",
000898 => x"E1A05000",
000899 => x"8A000098",
000900 => x"E3700004",
000901 => x"12844008",
000902 => x"1280600B",
000903 => x"0A000006",
000904 => x"EBFFFCE8",
000905 => x"E3700001",
000906 => x"0AFFFFFC",
000907 => x"E1560004",
000908 => x"E5C40000",
000909 => x"E2844001",
000910 => x"1AFFFFF8",
000911 => x"E59F02D0",
000912 => x"EBFFFDB9",
000913 => x"E59F02CC",
000914 => x"EBFFFDB7",
000915 => x"E375000C",
000916 => x"0A00000F",
000917 => x"E3A04000",
000918 => x"E285700C",
000919 => x"E1A06004",
000920 => x"E5D45000",
000921 => x"E3A00077",
000922 => x"E1A01008",
000923 => x"E1A02006",
000924 => x"E3A03002",
000925 => x"E58D5000",
000926 => x"EBFFFD14",
000927 => x"E3500000",
000928 => x"1AFFFFF7",
000929 => x"E2844001",
000930 => x"E1540007",
000931 => x"E1A06004",
000932 => x"1AFFFFF2",
000933 => x"E59F0280",
000934 => x"EBFFFDA3",
000935 => x"EAFFFFB6",
000936 => x"E1A00004",
000937 => x"EBFFFCCD",
000938 => x"E59F0270",
000939 => x"EBFFFD9E",
000940 => x"E59F026C",
000941 => x"EBFFFD9C",
000942 => x"E59F0268",
000943 => x"EBFFFD9A",
000944 => x"E59F0264",
000945 => x"EBFFFD98",
000946 => x"E59F0260",
000947 => x"EBFFFD96",
000948 => x"E59F025C",
000949 => x"EBFFFD94",
000950 => x"E59F0258",
000951 => x"EBFFFD92",
000952 => x"E59F0254",
000953 => x"EBFFFD90",
000954 => x"E59F0250",
000955 => x"EBFFFD8E",
000956 => x"E59F024C",
000957 => x"EBFFFD8C",
000958 => x"E59F0248",
000959 => x"EBFFFD8A",
000960 => x"E59F0244",
000961 => x"EBFFFD88",
000962 => x"E59F0240",
000963 => x"EBFFFD86",
000964 => x"E59F023C",
000965 => x"EBFFFD84",
000966 => x"E59F0238",
000967 => x"EBFFFD82",
000968 => x"E59F0234",
000969 => x"EBFFFD80",
000970 => x"E59F0230",
000971 => x"EBFFFD7E",
000972 => x"E59F022C",
000973 => x"EBFFFD7C",
000974 => x"E59F0228",
000975 => x"EBFFFD7A",
000976 => x"E59F0224",
000977 => x"EBFFFD78",
000978 => x"EAFFFE51",
000979 => x"E5DD3011",
000980 => x"E3530042",
000981 => x"1AFFFEEB",
000982 => x"E5DD3012",
000983 => x"E3530052",
000984 => x"1AFFFEE8",
000985 => x"E3A01004",
000986 => x"E3A02000",
000987 => x"E1A0000A",
000988 => x"EBFFFD7B",
000989 => x"E1A0000A",
000990 => x"EBFFFDFC",
000991 => x"E3A03C7F",
000992 => x"E28330F8",
000993 => x"E1500003",
000994 => x"8A000039",
000995 => x"E2804401",
000996 => x"E2844004",
000997 => x"E3540401",
000998 => x"0A000009",
000999 => x"E3A05401",
001000 => x"E3A01004",
001001 => x"E3A02000",
001002 => x"E1A0000A",
001003 => x"EBFFFD6C",
001004 => x"E1A0000A",
001005 => x"EBFFFDED",
001006 => x"E4850004",
001007 => x"E1550004",
001008 => x"1AFFFFF6",
001009 => x"EBFFFDF1",
001010 => x"EAFFFE31",
001011 => x"E1A00004",
001012 => x"EBFFFC82",
001013 => x"E59F0194",
001014 => x"EBFFFD53",
001015 => x"E1A0000A",
001016 => x"E3A01002",
001017 => x"E3A02001",
001018 => x"EBFFFD5D",
001019 => x"E1A0000A",
001020 => x"E3A01002",
001021 => x"EBFFFDC2",
001022 => x"E21060FF",
001023 => x"0AFFFE91",
001024 => x"E59F016C",
001025 => x"EBFFFD48",
001026 => x"E59F0168",
001027 => x"EBFFFD46",
001028 => x"EBFFFC6C",
001029 => x"E3700001",
001030 => x"0AFFFFFC",
001031 => x"EBFFFC69",
001032 => x"E3700001",
001033 => x"1AFFFFFC",
001034 => x"E3A05000",
001035 => x"EA000001",
001036 => x"E3540000",
001037 => x"AA000011",
001038 => x"E3A0C000",
001039 => x"E1A02005",
001040 => x"E1A01006",
001041 => x"E3A03002",
001042 => x"E3A00072",
001043 => x"E58DC000",
001044 => x"EBFFFC9E",
001045 => x"E1A04000",
001046 => x"EBFFFC5A",
001047 => x"E3700001",
001048 => x"E1A00004",
001049 => x"0AFFFFF1",
001050 => x"E59F010C",
001051 => x"EBFFFD2E",
001052 => x"EAFFFF23",
001053 => x"E59F0104",
001054 => x"EBFFFD2B",
001055 => x"EAFFFE04",
001056 => x"EBFFFC56",
001057 => x"E3A03801",
001058 => x"E2855001",
001059 => x"E2433001",
001060 => x"E1550003",
001061 => x"1AFFFFE7",
001062 => x"EAFFFF19",
001063 => x"000112C0",
001064 => x"0001130C",
001065 => x"00011354",
001066 => x"0001139C",
001067 => x"000113E4",
001068 => x"0001142C",
001069 => x"00011474",
001070 => x"000114E0",
001071 => x"00011518",
001072 => x"00011528",
001073 => x"000116B4",
001074 => x"00011718",
001075 => x"00011E1C",
001076 => x"00011658",
001077 => x"00011694",
001078 => x"00011744",
001079 => x"0001152C",
001080 => x"000115C4",
001081 => x"00011DA0",
001082 => x"00011DD0",
001083 => x"00011704",
001084 => x"00011DF8",
001085 => x"000115EC",
001086 => x"00011634",
001087 => x"000118F4",
001088 => x"00011928",
001089 => x"00011994",
001090 => x"00011764",
001091 => x"0001180C",
001092 => x"00011DEC",
001093 => x"000117C4",
001094 => x"000117DC",
001095 => x"000117FC",
001096 => x"000119D8",
001097 => x"000119F4",
001098 => x"00011A14",
001099 => x"00011A54",
001100 => x"00011A88",
001101 => x"00011AC4",
001102 => x"00011B00",
001103 => x"00011B24",
001104 => x"00011B60",
001105 => x"00011B7C",
001106 => x"00011B94",
001107 => x"00011BDC",
001108 => x"00011C1C",
001109 => x"00011C54",
001110 => x"00011C78",
001111 => x"00011CBC",
001112 => x"00011CFC",
001113 => x"00011D28",
001114 => x"00011D54",
001115 => x"00011D78",
001116 => x"00011830",
001117 => x"0001186C",
001118 => x"000118AC",
001119 => x"00011E40",
001120 => x"000115A0",
001121 => x"E10F3000",
001122 => x"E3C330C0",
001123 => x"E129F003",
001124 => x"E1A0F00E",
001125 => x"E10F3000",
001126 => x"E38330C0",
001127 => x"E129F003",
001128 => x"E1A0F00E",
001129 => x"00000000",
001130 => x"2030202D",
001131 => x"20626F6F",
001132 => x"74206672",
001133 => x"6F6D2063",
001134 => x"6F726520",
001135 => x"52414D20",
001136 => x"28737461",
001137 => x"72742061",
001138 => x"70706C69",
001139 => x"63617469",
001140 => x"6F6E290D",
001141 => x"0A203120",
001142 => x"2D207072",
001143 => x"6F677261",
001144 => x"6D20636F",
001145 => x"72652052",
001146 => x"414D2076",
001147 => x"69612055",
001148 => x"4152545F",
001149 => x"300D0A20",
001150 => x"32202D20",
001151 => x"636F7265",
001152 => x"2052414D",
001153 => x"2064756D",
001154 => x"700D0A00",
001155 => x"2033202D",
001156 => x"20626F6F",
001157 => x"74206672",
001158 => x"6F6D2049",
001159 => x"32432045",
001160 => x"4550524F",
001161 => x"4D0D0A20",
001162 => x"34202D20",
001163 => x"70726F67",
001164 => x"72616D20",
001165 => x"49324320",
001166 => x"45455052",
001167 => x"4F4D2076",
001168 => x"69612055",
001169 => x"4152545F",
001170 => x"300D0A20",
001171 => x"35202D20",
001172 => x"73686F77",
001173 => x"20636F6E",
001174 => x"74656E74",
001175 => x"206F6620",
001176 => x"49324320",
001177 => x"45455052",
001178 => x"4F4D0D0A",
001179 => x"00000000",
001180 => x"2061202D",
001181 => x"20617574",
001182 => x"6F6D6174",
001183 => x"69632062",
001184 => x"6F6F7420",
001185 => x"636F6E66",
001186 => x"69677572",
001187 => x"6174696F",
001188 => x"6E0D0A20",
001189 => x"68202D20",
001190 => x"68656C70",
001191 => x"0D0A2072",
001192 => x"202D2072",
001193 => x"65737461",
001194 => x"72742073",
001195 => x"79737465",
001196 => x"6D0D0A0D",
001197 => x"0A53656C",
001198 => x"6563743A",
001199 => x"20000000",
001200 => x"0D0A0D0A",
001201 => x"0D0A2B2D",
001202 => x"2D2D2D2D",
001203 => x"2D2D2D2D",
001204 => x"2D2D2D2D",
001205 => x"2D2D2D2D",
001206 => x"2D2D2D2D",
001207 => x"2D2D2D2D",
001208 => x"2D2D2D2D",
001209 => x"2D2D2D2D",
001210 => x"2D2D2D2D",
001211 => x"2D2D2D2D",
001212 => x"2D2D2D2D",
001213 => x"2D2D2D2D",
001214 => x"2D2D2D2D",
001215 => x"2D2D2D2D",
001216 => x"2D2D2D2D",
001217 => x"2D2D2D2B",
001218 => x"0D0A0000",
001219 => x"7C202020",
001220 => x"203C3C3C",
001221 => x"2053544F",
001222 => x"524D2043",
001223 => x"6F726520",
001224 => x"50726F63",
001225 => x"6573736F",
001226 => x"72205379",
001227 => x"7374656D",
001228 => x"202D2042",
001229 => x"79205374",
001230 => x"65706861",
001231 => x"6E204E6F",
001232 => x"6C74696E",
001233 => x"67203E3E",
001234 => x"3E202020",
001235 => x"207C0D0A",
001236 => x"00000000",
001237 => x"2B2D2D2D",
001238 => x"2D2D2D2D",
001239 => x"2D2D2D2D",
001240 => x"2D2D2D2D",
001241 => x"2D2D2D2D",
001242 => x"2D2D2D2D",
001243 => x"2D2D2D2D",
001244 => x"2D2D2D2D",
001245 => x"2D2D2D2D",
001246 => x"2D2D2D2D",
001247 => x"2D2D2D2D",
001248 => x"2D2D2D2D",
001249 => x"2D2D2D2D",
001250 => x"2D2D2D2D",
001251 => x"2D2D2D2D",
001252 => x"2D2D2D2D",
001253 => x"2D2B0D0A",
001254 => x"00000000",
001255 => x"7C202020",
001256 => x"20202020",
001257 => x"2020426F",
001258 => x"6F746C6F",
001259 => x"61646572",
001260 => x"20666F72",
001261 => x"2053544F",
001262 => x"524D2053",
001263 => x"6F432020",
001264 => x"20566572",
001265 => x"73696F6E",
001266 => x"3A203230",
001267 => x"31323035",
001268 => x"32342D44",
001269 => x"20202020",
001270 => x"20202020",
001271 => x"207C0D0A",
001272 => x"00000000",
001273 => x"7C202020",
001274 => x"20202020",
001275 => x"20202020",
001276 => x"20202020",
001277 => x"436F6E74",
001278 => x"6163743A",
001279 => x"2073746E",
001280 => x"6F6C7469",
001281 => x"6E674067",
001282 => x"6F6F676C",
001283 => x"656D6169",
001284 => x"6C2E636F",
001285 => x"6D202020",
001286 => x"20202020",
001287 => x"20202020",
001288 => x"20202020",
001289 => x"207C0D0A",
001290 => x"00000000",
001291 => x"2B2D2D2D",
001292 => x"2D2D2D2D",
001293 => x"2D2D2D2D",
001294 => x"2D2D2D2D",
001295 => x"2D2D2D2D",
001296 => x"2D2D2D2D",
001297 => x"2D2D2D2D",
001298 => x"2D2D2D2D",
001299 => x"2D2D2D2D",
001300 => x"2D2D2D2D",
001301 => x"2D2D2D2D",
001302 => x"2D2D2D2D",
001303 => x"2D2D2D2D",
001304 => x"2D2D2D2D",
001305 => x"2D2D2D2D",
001306 => x"2D2D2D2D",
001307 => x"2D2B0D0A",
001308 => x"0D0A0000",
001309 => x"203C2057",
001310 => x"656C636F",
001311 => x"6D652074",
001312 => x"6F207468",
001313 => x"65205354",
001314 => x"4F524D20",
001315 => x"536F4320",
001316 => x"626F6F74",
001317 => x"6C6F6164",
001318 => x"65722063",
001319 => x"6F6E736F",
001320 => x"6C652120",
001321 => x"3E0D0A20",
001322 => x"3C205365",
001323 => x"6C656374",
001324 => x"20616E20",
001325 => x"6F706572",
001326 => x"6174696F",
001327 => x"6E206672",
001328 => x"6F6D2074",
001329 => x"6865206D",
001330 => x"656E7520",
001331 => x"62656C6F",
001332 => x"77206F72",
001333 => x"20707265",
001334 => x"7373203E",
001335 => x"0D0A0000",
001336 => x"203C2074",
001337 => x"68652062",
001338 => x"6F6F7420",
001339 => x"6B657920",
001340 => x"666F7220",
001341 => x"696D6D65",
001342 => x"64696174",
001343 => x"65206170",
001344 => x"706C6963",
001345 => x"6174696F",
001346 => x"6E207374",
001347 => x"6172742E",
001348 => x"203E0D0A",
001349 => x"0D0A0000",
001350 => x"204C6F61",
001351 => x"64204164",
001352 => x"64726573",
001353 => x"733A2000",
001354 => x"0A0D0000",
001355 => x"0D0A0D0A",
001356 => x"4170706C",
001357 => x"69636174",
001358 => x"696F6E20",
001359 => x"77696C6C",
001360 => x"20737461",
001361 => x"72742061",
001362 => x"75746F6D",
001363 => x"61746963",
001364 => x"616C6C79",
001365 => x"20616674",
001366 => x"65722064",
001367 => x"6F776E6C",
001368 => x"6F61642E",
001369 => x"0D0A2D3E",
001370 => x"20576169",
001371 => x"74696E67",
001372 => x"20666F72",
001373 => x"20277374",
001374 => x"6F726D5F",
001375 => x"70726F67",
001376 => x"72616D2E",
001377 => x"62696E27",
001378 => x"20696E20",
001379 => x"62797465",
001380 => x"2D737472",
001381 => x"65616D20",
001382 => x"6D6F6465",
001383 => x"2E2E2E00",
001384 => x"20455252",
001385 => x"4F522120",
001386 => x"50726F67",
001387 => x"72616D20",
001388 => x"66696C65",
001389 => x"20746F6F",
001390 => x"20626967",
001391 => x"210D0A0D",
001392 => x"0A000000",
001393 => x"20496E76",
001394 => x"616C6964",
001395 => x"2070726F",
001396 => x"6772616D",
001397 => x"6D696E67",
001398 => x"2066696C",
001399 => x"65210D0A",
001400 => x"0D0A5365",
001401 => x"6C656374",
001402 => x"3A200000",
001403 => x"0D0A0D0A",
001404 => x"41626F72",
001405 => x"74206475",
001406 => x"6D70696E",
001407 => x"67206279",
001408 => x"20707265",
001409 => x"7373696E",
001410 => x"6720616E",
001411 => x"79206B65",
001412 => x"792E0D0A",
001413 => x"50726573",
001414 => x"7320616E",
001415 => x"79206B65",
001416 => x"7920746F",
001417 => x"20636F6E",
001418 => x"74696E75",
001419 => x"652E0D0A",
001420 => x"0D0A0000",
001421 => x"0D0A0D0A",
001422 => x"44756D70",
001423 => x"696E6720",
001424 => x"636F6D70",
001425 => x"6C657465",
001426 => x"642E0D0A",
001427 => x"0D0A5365",
001428 => x"6C656374",
001429 => x"3A200000",
001430 => x"0D0A0D0A",
001431 => x"456E7465",
001432 => x"72206465",
001433 => x"76696365",
001434 => x"20616464",
001435 => x"72657373",
001436 => x"20283278",
001437 => x"20686578",
001438 => x"5F636861",
001439 => x"72732C20",
001440 => x"73657420",
001441 => x"4C534220",
001442 => x"746F2027",
001443 => x"3027293A",
001444 => x"20000000",
001445 => x"20496E76",
001446 => x"616C6964",
001447 => x"20616464",
001448 => x"72657373",
001449 => x"210D0A0D",
001450 => x"0A53656C",
001451 => x"6563743A",
001452 => x"20000000",
001453 => x"0D0A4170",
001454 => x"706C6963",
001455 => x"6174696F",
001456 => x"6E207769",
001457 => x"6C6C2073",
001458 => x"74617274",
001459 => x"20617574",
001460 => x"6F6D6174",
001461 => x"6963616C",
001462 => x"6C792061",
001463 => x"66746572",
001464 => x"2075706C",
001465 => x"6F61642E",
001466 => x"0D0A2D3E",
001467 => x"204C6F61",
001468 => x"64696E67",
001469 => x"20626F6F",
001470 => x"7420696D",
001471 => x"6167652E",
001472 => x"2E2E0000",
001473 => x"2055706C",
001474 => x"6F616420",
001475 => x"636F6D70",
001476 => x"6C657465",
001477 => x"0D0A0000",
001478 => x"20496E76",
001479 => x"616C6964",
001480 => x"20626F6F",
001481 => x"74206465",
001482 => x"76696365",
001483 => x"206F7220",
001484 => x"66696C65",
001485 => x"210D0A0D",
001486 => x"0A53656C",
001487 => x"6563743A",
001488 => x"20000000",
001489 => x"0D0A496E",
001490 => x"76616C69",
001491 => x"64206164",
001492 => x"64726573",
001493 => x"73210D0A",
001494 => x"0D0A5365",
001495 => x"6C656374",
001496 => x"3A200000",
001497 => x"0D0A4461",
001498 => x"74612077",
001499 => x"696C6C20",
001500 => x"6F766572",
001501 => x"77726974",
001502 => x"65205241",
001503 => x"4D20636F",
001504 => x"6E74656E",
001505 => x"74210D0A",
001506 => x"2D3E2057",
001507 => x"61697469",
001508 => x"6E672066",
001509 => x"6F722027",
001510 => x"73746F72",
001511 => x"6D5F7072",
001512 => x"6F677261",
001513 => x"6D2E6269",
001514 => x"6E272069",
001515 => x"6E206279",
001516 => x"74652D73",
001517 => x"74726561",
001518 => x"6D206D6F",
001519 => x"64652E2E",
001520 => x"2E000000",
001521 => x"20446F77",
001522 => x"6E6C6F61",
001523 => x"6420636F",
001524 => x"6D706C65",
001525 => x"7465640D",
001526 => x"0A000000",
001527 => x"57726974",
001528 => x"696E6720",
001529 => x"62756666",
001530 => x"65722074",
001531 => x"6F206932",
001532 => x"63204545",
001533 => x"50524F4D",
001534 => x"2E2E2E00",
001535 => x"20436F6D",
001536 => x"706C6574",
001537 => x"65640D0A",
001538 => x"0D0A0000",
001539 => x"20496E76",
001540 => x"616C6964",
001541 => x"20626F6F",
001542 => x"74206465",
001543 => x"76696365",
001544 => x"206F7220",
001545 => x"66696C65",
001546 => x"210D0A0D",
001547 => x"0A000000",
001548 => x"0D0A0D0A",
001549 => x"456E7465",
001550 => x"72206465",
001551 => x"76696365",
001552 => x"20616464",
001553 => x"72657373",
001554 => x"20283220",
001555 => x"6865782D",
001556 => x"63686172",
001557 => x"732C2073",
001558 => x"6574204C",
001559 => x"53422074",
001560 => x"6F202730",
001561 => x"27293A20",
001562 => x"00000000",
001563 => x"0D0A0D0A",
001564 => x"41626F72",
001565 => x"74206475",
001566 => x"6D70696E",
001567 => x"67206279",
001568 => x"20707265",
001569 => x"7373696E",
001570 => x"6720616E",
001571 => x"79206B65",
001572 => x"792E2049",
001573 => x"66206E6F",
001574 => x"20646174",
001575 => x"61206973",
001576 => x"2073686F",
001577 => x"776E2C0D",
001578 => x"0A000000",
001579 => x"74686520",
001580 => x"73656C65",
001581 => x"63746564",
001582 => x"20646576",
001583 => x"69636520",
001584 => x"6973206E",
001585 => x"6F742072",
001586 => x"6573706F",
001587 => x"6E64696E",
001588 => x"672E2050",
001589 => x"72657373",
001590 => x"20616E79",
001591 => x"206B6579",
001592 => x"20746F20",
001593 => x"636F6E74",
001594 => x"696E7565",
001595 => x"2E0D0A0D",
001596 => x"0A000000",
001597 => x"0D0A0D0A",
001598 => x"4175746F",
001599 => x"6D617469",
001600 => x"6320626F",
001601 => x"6F742063",
001602 => x"6F6E6669",
001603 => x"67757261",
001604 => x"74696F6E",
001605 => x"20666F72",
001606 => x"20706F77",
001607 => x"65722D75",
001608 => x"703A0D0A",
001609 => x"00000000",
001610 => x"5B333231",
001611 => x"305D2063",
001612 => x"6F6E6669",
001613 => x"67757261",
001614 => x"74696F6E",
001615 => x"20444950",
001616 => x"20737769",
001617 => x"7463680D",
001618 => x"0A203030",
001619 => x"3030202D",
001620 => x"20537461",
001621 => x"72742062",
001622 => x"6F6F746C",
001623 => x"6F616465",
001624 => x"7220636F",
001625 => x"6E736F6C",
001626 => x"650D0A20",
001627 => x"30303031",
001628 => x"202D2041",
001629 => x"75746F6D",
001630 => x"61746963",
001631 => x"20626F6F",
001632 => x"74206672",
001633 => x"6F6D2063",
001634 => x"6F726520",
001635 => x"52414D0D",
001636 => x"0A000000",
001637 => x"20303031",
001638 => x"30202D20",
001639 => x"4175746F",
001640 => x"6D617469",
001641 => x"6320626F",
001642 => x"6F742066",
001643 => x"726F6D20",
001644 => x"49324320",
001645 => x"45455052",
001646 => x"4F4D2028",
001647 => x"41646472",
001648 => x"65737320",
001649 => x"30784130",
001650 => x"290D0A0D",
001651 => x"0A53656C",
001652 => x"6563743A",
001653 => x"20000000",
001654 => x"0D0A0D0A",
001655 => x"53544F52",
001656 => x"4D20536F",
001657 => x"4320626F",
001658 => x"6F746C6F",
001659 => x"61646572",
001660 => x"0D0A0000",
001661 => x"2730273A",
001662 => x"20457865",
001663 => x"63757465",
001664 => x"2070726F",
001665 => x"6772616D",
001666 => x"20696E20",
001667 => x"52414D2E",
001668 => x"0D0A0000",
001669 => x"2731273A",
001670 => x"20577269",
001671 => x"74652027",
001672 => x"73746F72",
001673 => x"6D5F7072",
001674 => x"6F677261",
001675 => x"6D2E6269",
001676 => x"6E272074",
001677 => x"6F207468",
001678 => x"6520636F",
001679 => x"72652773",
001680 => x"2052414D",
001681 => x"20766961",
001682 => x"20554152",
001683 => x"542E0D0A",
001684 => x"00000000",
001685 => x"2732273A",
001686 => x"20507269",
001687 => x"6E742063",
001688 => x"75727265",
001689 => x"6E742063",
001690 => x"6F6E7465",
001691 => x"6E74206F",
001692 => x"6620636F",
001693 => x"6D706C65",
001694 => x"74652063",
001695 => x"6F726520",
001696 => x"52414D2E",
001697 => x"0D0A0000",
001698 => x"2733273A",
001699 => x"204C6F61",
001700 => x"6420626F",
001701 => x"6F742069",
001702 => x"6D616765",
001703 => x"2066726F",
001704 => x"6D204545",
001705 => x"50524F4D",
001706 => x"20616E64",
001707 => x"20737461",
001708 => x"72742061",
001709 => x"70706C69",
001710 => x"63617469",
001711 => x"6F6E2E0D",
001712 => x"0A000000",
001713 => x"2734273A",
001714 => x"20577269",
001715 => x"74652027",
001716 => x"73746F72",
001717 => x"6D5F7072",
001718 => x"6F677261",
001719 => x"6D2E6269",
001720 => x"6E272074",
001721 => x"6F204932",
001722 => x"43204545",
001723 => x"50524F4D",
001724 => x"20766961",
001725 => x"20554152",
001726 => x"542E0D0A",
001727 => x"00000000",
001728 => x"2735273A",
001729 => x"20507269",
001730 => x"6E742063",
001731 => x"6F6E7465",
001732 => x"6E74206F",
001733 => x"66204932",
001734 => x"43204545",
001735 => x"50524F4D",
001736 => x"2E0D0A00",
001737 => x"2761273A",
001738 => x"2053686F",
001739 => x"77204449",
001740 => x"50207377",
001741 => x"69746368",
001742 => x"20636F6E",
001743 => x"66696775",
001744 => x"72617469",
001745 => x"6F6E7320",
001746 => x"666F7220",
001747 => x"6175746F",
001748 => x"6D617469",
001749 => x"6320626F",
001750 => x"6F742E0D",
001751 => x"0A000000",
001752 => x"2768273A",
001753 => x"2053686F",
001754 => x"77207468",
001755 => x"69732073",
001756 => x"63726565",
001757 => x"6E2E0D0A",
001758 => x"00000000",
001759 => x"2772273A",
001760 => x"20526573",
001761 => x"65742073",
001762 => x"79737465",
001763 => x"6D2E0D0A",
001764 => x"0D0A0000",
001765 => x"426F6F74",
001766 => x"20454550",
001767 => x"524F4D3A",
001768 => x"20323478",
001769 => x"786E6E6E",
001770 => x"20286C69",
001771 => x"6B652032",
001772 => x"34414136",
001773 => x"34292C20",
001774 => x"37206269",
001775 => x"74206164",
001776 => x"64726573",
001777 => x"73202B20",
001778 => x"646F6E74",
001779 => x"2D636172",
001780 => x"65206269",
001781 => x"742C0D0A",
001782 => x"00000000",
001783 => x"636F6E6E",
001784 => x"65637465",
001785 => x"6420746F",
001786 => x"20493243",
001787 => x"5F434F4E",
001788 => x"54524F4C",
001789 => x"4C45525F",
001790 => x"302C206F",
001791 => x"70657261",
001792 => x"74696E67",
001793 => x"20667265",
001794 => x"7175656E",
001795 => x"63792069",
001796 => x"73203130",
001797 => x"306B487A",
001798 => x"2C0D0A00",
001799 => x"6D617869",
001800 => x"6D756D20",
001801 => x"45455052",
001802 => x"4F4D2073",
001803 => x"697A6520",
001804 => x"3D203635",
001805 => x"35333620",
001806 => x"62797465",
001807 => x"203D3E20",
001808 => x"31362062",
001809 => x"69742061",
001810 => x"64647265",
001811 => x"73736573",
001812 => x"2C0D0A00",
001813 => x"66697865",
001814 => x"6420626F",
001815 => x"6F742064",
001816 => x"65766963",
001817 => x"65206164",
001818 => x"64726573",
001819 => x"733A2030",
001820 => x"7841300D",
001821 => x"0A0D0A00",
001822 => x"5465726D",
001823 => x"696E616C",
001824 => x"20736574",
001825 => x"75703A20",
001826 => x"39363030",
001827 => x"20626175",
001828 => x"642C2038",
001829 => x"20646174",
001830 => x"61206269",
001831 => x"74732C20",
001832 => x"6E6F2070",
001833 => x"61726974",
001834 => x"792C2031",
001835 => x"2073746F",
001836 => x"70206269",
001837 => x"740D0A0D",
001838 => x"0A000000",
001839 => x"466F7220",
001840 => x"6D6F7265",
001841 => x"20696E66",
001842 => x"6F726D61",
001843 => x"74696F6E",
001844 => x"20736565",
001845 => x"20746865",
001846 => x"2053544F",
001847 => x"524D2043",
001848 => x"6F726520",
001849 => x"2F205354",
001850 => x"4F524D20",
001851 => x"536F4320",
001852 => x"64617461",
001853 => x"73686565",
001854 => x"740D0A00",
001855 => x"68747470",
001856 => x"3A2F2F6F",
001857 => x"70656E63",
001858 => x"6F726573",
001859 => x"2E6F7267",
001860 => x"2F70726F",
001861 => x"6A656374",
001862 => x"2C73746F",
001863 => x"726D5F63",
001864 => x"6F72650D",
001865 => x"0A000000",
001866 => x"68747470",
001867 => x"3A2F2F6F",
001868 => x"70656E63",
001869 => x"6F726573",
001870 => x"2E6F7267",
001871 => x"2F70726F",
001872 => x"6A656374",
001873 => x"2C73746F",
001874 => x"726D5F73",
001875 => x"6F630D0A",
001876 => x"00000000",
001877 => x"436F6E74",
001878 => x"6163743A",
001879 => x"2073746E",
001880 => x"6F6C7469",
001881 => x"6E674067",
001882 => x"6F6F676C",
001883 => x"656D6169",
001884 => x"6C2E636F",
001885 => x"6D0D0A00",
001886 => x"28632920",
001887 => x"32303132",
001888 => x"20627920",
001889 => x"53746570",
001890 => x"68616E20",
001891 => x"4E6F6C74",
001892 => x"696E670D",
001893 => x"0A0D0A53",
001894 => x"656C6563",
001895 => x"743A2000",
001896 => x"0D0A0D0A",
001897 => x"5765276C",
001898 => x"6C207365",
001899 => x"6E642079",
001900 => x"6F752062",
001901 => x"61636B20",
001902 => x"2D20746F",
001903 => x"20746865",
001904 => x"20667574",
001905 => x"75726521",
001906 => x"2E0D0A0D",
001907 => x"0A000000",
001908 => x"202D2044",
001909 => x"6F63746F",
001910 => x"7220456D",
001911 => x"6D657420",
001912 => x"4C2E2042",
001913 => x"726F776E",
001914 => x"0D0A0D0A",
001915 => x"53656C65",
001916 => x"63743A20",
001917 => x"00000000",
001918 => x"20496E76",
001919 => x"616C6964",
001920 => x"206F7065",
001921 => x"72617469",
001922 => x"6F6E210D",
001923 => x"0A547279",
001924 => x"20616761",
001925 => x"696E3A20",
001926 => x"00000000",
001927 => x"0D0A0D0A",
001928 => x"2D3E2053",
001929 => x"74617274",
001930 => x"696E6720",
001931 => x"6170706C",
001932 => x"69636174",
001933 => x"696F6E2E",
001934 => x"2E2E0D0A",
001935 => x"0D0A0000",
001936 => x"0D0A0D0A",
001937 => x"41626F72",
001938 => x"74656421",
001939 => x"00000000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;