-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
	--bootloader_sdram
000000 => x"EA000006",
000001 => x"EAFFFFFE",
000002 => x"EAFFFFFE",
000003 => x"EAFFFFFE",
000004 => x"EAFFFFFE",
000005 => x"E1A00000",
000006 => x"EAFFFFFE",
000007 => x"EAFFFFFE",
000008 => x"E59F0040",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA018",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"E1A04000",
000023 => x"E3A00000",
000024 => x"E1A0F004",
000025 => x"EAFFFFFE",
000026 => x"00002000",
000027 => x"000107BC",
000028 => x"E3E03A0F",
000029 => x"E5131FFB",
000030 => x"E20020FF",
000031 => x"E3A00001",
000032 => x"E0010210",
000033 => x"E1A0F00E",
000034 => x"E3E03A0F",
000035 => x"E5130FFB",
000036 => x"E1A0F00E",
000037 => x"E3E01A0F",
000038 => x"E5113FFF",
000039 => x"E20000FF",
000040 => x"E3A02001",
000041 => x"E1833012",
000042 => x"E5013FFF",
000043 => x"E1A0F00E",
000044 => x"E20000FF",
000045 => x"E3A02001",
000046 => x"E1A02012",
000047 => x"E3E01A0F",
000048 => x"E5113FFF",
000049 => x"E1E02002",
000050 => x"E0033002",
000051 => x"E5013FFF",
000052 => x"E1A0F00E",
000053 => x"E3E01A0F",
000054 => x"E5113FFF",
000055 => x"E20000FF",
000056 => x"E3A02001",
000057 => x"E0233012",
000058 => x"E5013FFF",
000059 => x"E1A0F00E",
000060 => x"E3E03A0F",
000061 => x"E5030FFF",
000062 => x"E1A0F00E",
000063 => x"E20000FF",
000064 => x"E3500007",
000065 => x"E92D4010",
000066 => x"E3A0C000",
000067 => x"E3E0E0FF",
000068 => x"E20110FF",
000069 => x"8A000011",
000070 => x"E2403004",
000071 => x"E20330FF",
000072 => x"E3500003",
000073 => x"E1A0E183",
000074 => x"E3E04A0F",
000075 => x"E1A0C180",
000076 => x"9A000007",
000077 => x"E3A030FF",
000078 => x"E1A03E13",
000079 => x"E5142F8B",
000080 => x"E1E03003",
000081 => x"E0022003",
000082 => x"E1822E11",
000083 => x"E5042F8B",
000084 => x"E8BD8010",
000085 => x"E3A030FF",
000086 => x"E1A03C13",
000087 => x"E1E0E003",
000088 => x"E3E02A0F",
000089 => x"E5123F8F",
000090 => x"E003300E",
000091 => x"E1833C11",
000092 => x"E5023F8F",
000093 => x"E8BD8010",
000094 => x"E20000FF",
000095 => x"E3500007",
000096 => x"E3A02000",
000097 => x"8A00000A",
000098 => x"E2403004",
000099 => x"E3500003",
000100 => x"E20320FF",
000101 => x"9A000005",
000102 => x"E3E03A0F",
000103 => x"E5130F8B",
000104 => x"E1A02182",
000105 => x"E1A00230",
000106 => x"E20000FF",
000107 => x"E1A0F00E",
000108 => x"E1A02180",
000109 => x"E3E03A0F",
000110 => x"E5130F8F",
000111 => x"E1A00230",
000112 => x"E20000FF",
000113 => x"E1A0F00E",
000114 => x"E3E02A0F",
000115 => x"E5123EFB",
000116 => x"E3130002",
000117 => x"E3E00000",
000118 => x"15120EFF",
000119 => x"E1A0F00E",
000120 => x"E3E02A0F",
000121 => x"E5123EFB",
000122 => x"E3130001",
000123 => x"0AFFFFFC",
000124 => x"E20030FF",
000125 => x"E5023EFF",
000126 => x"E1A0F00E",
000127 => x"E20000FF",
000128 => x"E3500001",
000129 => x"E3812B01",
000130 => x"03E03A0F",
000131 => x"E3811B09",
000132 => x"13E03A0F",
000133 => x"05031CFF",
000134 => x"15032CFF",
000135 => x"E1A0F00E",
000136 => x"E3E03A0F",
000137 => x"E5030CFB",
000138 => x"E1A0F00E",
000139 => x"E3E02A0F",
000140 => x"E5123CFF",
000141 => x"E3130C01",
000142 => x"1AFFFFFC",
000143 => x"E5020CEF",
000144 => x"E5123CFF",
000145 => x"E3833C01",
000146 => x"E5023CFF",
000147 => x"E3E02A0F",
000148 => x"E5123CFF",
000149 => x"E3130C01",
000150 => x"1AFFFFFC",
000151 => x"E5120CEF",
000152 => x"E1A0F00E",
000153 => x"E3E01A0F",
000154 => x"E5113CF7",
000155 => x"E20000FF",
000156 => x"E3A02001",
000157 => x"E1833012",
000158 => x"E5013CF7",
000159 => x"E1A0F00E",
000160 => x"E20000FF",
000161 => x"E3A02001",
000162 => x"E1A02012",
000163 => x"E3E01A0F",
000164 => x"E5113CF7",
000165 => x"E1E02002",
000166 => x"E0033002",
000167 => x"E5013CF7",
000168 => x"E1A0F00E",
000169 => x"E3E02A0F",
000170 => x"E5123BE7",
000171 => x"E1A01420",
000172 => x"E3C33080",
000173 => x"E5023BE7",
000174 => x"E5020BEF",
000175 => x"E5021BEB",
000176 => x"E5123BE7",
000177 => x"E3833080",
000178 => x"E5023BE7",
000179 => x"E1A0F00E",
000180 => x"E92D4030",
000181 => x"E3A0C090",
000182 => x"E20140FE",
000183 => x"E3E0EA0F",
000184 => x"E5DD500F",
000185 => x"E20000FF",
000186 => x"E50E4BE3",
000187 => x"E20110FF",
000188 => x"E50ECBFF",
000189 => x"E1A04002",
000190 => x"E203C0FF",
000191 => x"E51E3BFF",
000192 => x"E3130002",
000193 => x"1AFFFFFC",
000194 => x"E51E3BFF",
000195 => x"E3130080",
000196 => x"13E00000",
000197 => x"18BD8030",
000198 => x"E35C0000",
000199 => x"0A000012",
000200 => x"E24C3001",
000201 => x"E203C0FF",
000202 => x"E35C0001",
000203 => x"01A02424",
000204 => x"03E03A0F",
000205 => x"13E03A0F",
000206 => x"05032BE3",
000207 => x"15034BE3",
000208 => x"E3E02A0F",
000209 => x"E3A03010",
000210 => x"E5023BFF",
000211 => x"E5123BFF",
000212 => x"E3130002",
000213 => x"1AFFFFFC",
000214 => x"E5123BFF",
000215 => x"E3130080",
000216 => x"0AFFFFEC",
000217 => x"E3E00001",
000218 => x"E8BD8030",
000219 => x"E3500077",
000220 => x"1A00000C",
000221 => x"E3E03A0F",
000222 => x"E3A02050",
000223 => x"E5035BE3",
000224 => x"E5032BFF",
000225 => x"E1A02003",
000226 => x"E5123BFF",
000227 => x"E3130002",
000228 => x"1AFFFFFC",
000229 => x"E5123BFF",
000230 => x"E2130080",
000231 => x"08BD8030",
000232 => x"E3E00002",
000233 => x"E8BD8030",
000234 => x"E3500072",
000235 => x"13E00003",
000236 => x"18BD8030",
000237 => x"E3813001",
000238 => x"E3E02A0F",
000239 => x"E3A01090",
000240 => x"E5023BE3",
000241 => x"E5021BFF",
000242 => x"E5123BFF",
000243 => x"E3130002",
000244 => x"1AFFFFFC",
000245 => x"E5123BFF",
000246 => x"E3130080",
000247 => x"1AFFFFEF",
000248 => x"E3A03068",
000249 => x"E5023BFF",
000250 => x"E3E00A0F",
000251 => x"E5103BFF",
000252 => x"E3130002",
000253 => x"1AFFFFFC",
000254 => x"E5100BE3",
000255 => x"E8BD8030",
000256 => x"E20000FF",
000257 => x"E350000F",
000258 => x"979FF100",
000259 => x"EA00000F",
000260 => x"000104D0",
000261 => x"000104C8",
000262 => x"000104C0",
000263 => x"000104B8",
000264 => x"000104B0",
000265 => x"000104A8",
000266 => x"000104A0",
000267 => x"00010498",
000268 => x"00010490",
000269 => x"00010488",
000270 => x"00010480",
000271 => x"00010478",
000272 => x"00010470",
000273 => x"00010468",
000274 => x"00010460",
000275 => x"00010458",
000276 => x"E3A00000",
000277 => x"E1A0F00E",
000278 => x"EE1F0F1F",
000279 => x"E1A0F00E",
000280 => x"EE1E0F1E",
000281 => x"E1A0F00E",
000282 => x"EE1D0F1D",
000283 => x"E1A0F00E",
000284 => x"EE1C0F1C",
000285 => x"E1A0F00E",
000286 => x"EE1B0F1B",
000287 => x"E1A0F00E",
000288 => x"EE1A0F1A",
000289 => x"E1A0F00E",
000290 => x"EE190F19",
000291 => x"E1A0F00E",
000292 => x"EE180F18",
000293 => x"E1A0F00E",
000294 => x"EE170F17",
000295 => x"E1A0F00E",
000296 => x"EE160F16",
000297 => x"E1A0F00E",
000298 => x"EE150F15",
000299 => x"E1A0F00E",
000300 => x"EE140F14",
000301 => x"E1A0F00E",
000302 => x"EE130F13",
000303 => x"E1A0F00E",
000304 => x"EE120F12",
000305 => x"E1A0F00E",
000306 => x"EE110F11",
000307 => x"E1A0F00E",
000308 => x"EE100F10",
000309 => x"E1A0F00E",
000310 => x"E20110FF",
000311 => x"E2411006",
000312 => x"E3510007",
000313 => x"979FF101",
000314 => x"EA000008",
000315 => x"00010514",
000316 => x"00010510",
000317 => x"00010510",
000318 => x"00010510",
000319 => x"00010510",
000320 => x"0001051C",
000321 => x"00010524",
000322 => x"0001050C",
000323 => x"EE0D0F1D",
000324 => x"E1A0F00E",
000325 => x"EE060F16",
000326 => x"E1A0F00E",
000327 => x"EE0B0F1B",
000328 => x"E1A0F00E",
000329 => x"EE0C0F1C",
000330 => x"E1A0F00E",
000331 => x"E92D4010",
000332 => x"E1A04000",
000333 => x"E5D00000",
000334 => x"E3500000",
000335 => x"1A000003",
000336 => x"EA000005",
000337 => x"E5F40001",
000338 => x"E3500000",
000339 => x"0A000002",
000340 => x"EBFFFF22",
000341 => x"E3500000",
000342 => x"CAFFFFF9",
000343 => x"E1A00004",
000344 => x"E8BD8010",
000345 => x"E92D4070",
000346 => x"E2514000",
000347 => x"E1A05000",
000348 => x"E20260FF",
000349 => x"DA00000B",
000350 => x"EBFFFF12",
000351 => x"E3700001",
000352 => x"E20030FF",
000353 => x"0A000005",
000354 => x"E3560001",
000355 => x"E5C53000",
000356 => x"E1A00003",
000357 => x"E2855001",
000358 => x"0A000005",
000359 => x"E2444001",
000360 => x"E3540000",
000361 => x"CAFFFFF3",
000362 => x"E59F300C",
000363 => x"E5C53000",
000364 => x"E8BD8070",
000365 => x"EBFFFF09",
000366 => x"EAFFFFF7",
000367 => x"00011190",
000368 => x"E92D4030",
000369 => x"E2514000",
000370 => x"E1A05000",
000371 => x"D8BD8030",
000372 => x"E4D50001",
000373 => x"EBFFFF01",
000374 => x"E2544001",
000375 => x"1AFFFFFB",
000376 => x"E8BD8030",
000377 => x"E92D4010",
000378 => x"E20240FF",
000379 => x"E3540008",
000380 => x"83A04008",
000381 => x"8A000001",
000382 => x"E3540000",
000383 => x"03A04001",
000384 => x"E1A02001",
000385 => x"E1A0E004",
000386 => x"E1A0310E",
000387 => x"E35E0001",
000388 => x"E2433004",
000389 => x"E1A0C000",
000390 => x"81A0C330",
000391 => x"E24E3001",
000392 => x"E20CC00F",
000393 => x"E203E0FF",
000394 => x"E35C0009",
000395 => x"E28C3030",
000396 => x"828C3037",
000397 => x"E35E0000",
000398 => x"E4C23001",
000399 => x"1AFFFFF1",
000400 => x"E2443001",
000401 => x"E20330FF",
000402 => x"E0813003",
000403 => x"E5C3E001",
000404 => x"E8BD8010",
000405 => x"E92D4010",
000406 => x"E1A04000",
000407 => x"E3540007",
000408 => x"E3A01010",
000409 => x"E3A00001",
000410 => x"9A000001",
000411 => x"E3A00000",
000412 => x"E8BD8010",
000413 => x"EBFFFEE0",
000414 => x"E3A00006",
000415 => x"EBFFFEF8",
000416 => x"E3A00000",
000417 => x"EBFFFEE8",
000418 => x"E1A00584",
000419 => x"E8BD4010",
000420 => x"EAFFFEE5",
000421 => x"E0603280",
000422 => x"E0800103",
000423 => x"E0800100",
000424 => x"E1A00200",
000425 => x"E3500000",
000426 => x"D1A0F00E",
000427 => x"E1A00000",
000428 => x"E2500001",
000429 => x"1AFFFFFC",
000430 => x"E1A0F00E",
000431 => x"E212C0FF",
000432 => x"0A00000B",
000433 => x"E5D02000",
000434 => x"E5D13000",
000435 => x"E1520003",
000436 => x"0A000004",
000437 => x"EA000008",
000438 => x"E5F02001",
000439 => x"E5F13001",
000440 => x"E1520003",
000441 => x"1A000004",
000442 => x"E24C3001",
000443 => x"E213C0FF",
000444 => x"1AFFFFF8",
000445 => x"E3A00001",
000446 => x"E1A0F00E",
000447 => x"E3A00000",
000448 => x"E1A0F00E",
000449 => x"E92D4030",
000450 => x"E1A04081",
000451 => x"E3540000",
000452 => x"E1A05000",
000453 => x"D3A00000",
000454 => x"D8BD8030",
000455 => x"E3A00000",
000456 => x"E1A01000",
000457 => x"E7D12005",
000458 => x"E2423030",
000459 => x"E082C200",
000460 => x"E3530009",
000461 => x"E242E041",
000462 => x"924C0030",
000463 => x"9A000007",
000464 => x"E0823200",
000465 => x"E35E0005",
000466 => x"E242C061",
000467 => x"92430037",
000468 => x"9A000002",
000469 => x"E0823200",
000470 => x"E35C0005",
000471 => x"92430057",
000472 => x"E2811001",
000473 => x"E1510004",
000474 => x"1AFFFFED",
000475 => x"E8BD8030",
000476 => x"E5D03003",
000477 => x"E5D02002",
000478 => x"E5D01000",
000479 => x"E1833402",
000480 => x"E5D00001",
000481 => x"E1833C01",
000482 => x"E1830800",
000483 => x"E1A0F00E",
000484 => x"E52DE004",
000485 => x"E59F0014",
000486 => x"EBFFFF63",
000487 => x"E59F0010",
000488 => x"EBFFFF61",
000489 => x"E59F000C",
000490 => x"E49DE004",
000491 => x"EAFFFF5E",
000492 => x"00011194",
000493 => x"000111F8",
000494 => x"0001125C",
000495 => x"E92D47F0",
000496 => x"E3A00000",
000497 => x"E24DD014",
000498 => x"EBFFFE48",
000499 => x"E3A0100D",
000500 => x"E3A000C3",
000501 => x"EBFFFF3F",
000502 => x"E3A00063",
000503 => x"EBFFFEB0",
000504 => x"E3A00006",
000505 => x"EBFFFF05",
000506 => x"E3A01006",
000507 => x"E3800008",
000508 => x"EBFFFF38",
000509 => x"E3A0000D",
000510 => x"EBFFFF00",
000511 => x"E1A008A0",
000512 => x"E1E00000",
000513 => x"E200000F",
000514 => x"E3500001",
000515 => x"03A04030",
000516 => x"028DA006",
000517 => x"028D900F",
000518 => x"0A000020",
000519 => x"E3500002",
000520 => x"0A00007E",
000521 => x"E59F085C",
000522 => x"EBFFFF3F",
000523 => x"E59F0858",
000524 => x"EBFFFF3D",
000525 => x"E59F0854",
000526 => x"EBFFFF3B",
000527 => x"E59F0850",
000528 => x"EBFFFF39",
000529 => x"E59F084C",
000530 => x"EBFFFF37",
000531 => x"E59F0848",
000532 => x"EBFFFF35",
000533 => x"E59F0844",
000534 => x"EBFFFF33",
000535 => x"E59F0840",
000536 => x"EBFFFF31",
000537 => x"E28DA006",
000538 => x"E59F0838",
000539 => x"EBFFFF2E",
000540 => x"E1A0100A",
000541 => x"E3A02008",
000542 => x"E3A00301",
000543 => x"EBFFFF58",
000544 => x"E1A0000A",
000545 => x"EBFFFF28",
000546 => x"E59F081C",
000547 => x"EBFFFF26",
000548 => x"EBFFFFBE",
000549 => x"E28D900F",
000550 => x"EBFFFE4A",
000551 => x"E1A04000",
000552 => x"E3A0000D",
000553 => x"EBFFFED5",
000554 => x"E3100801",
000555 => x"03A06001",
000556 => x"03A050A0",
000557 => x"1A00003D",
000558 => x"E3A04000",
000559 => x"E59F07EC",
000560 => x"EBFFFF19",
000561 => x"E1A01005",
000562 => x"E1A02004",
000563 => x"E3A03002",
000564 => x"E3A00072",
000565 => x"E58D4000",
000566 => x"EBFFFE7C",
000567 => x"E1A01005",
000568 => x"E5CD000F",
000569 => x"E3A02001",
000570 => x"E3A03002",
000571 => x"E3A00072",
000572 => x"E58D4000",
000573 => x"EBFFFE75",
000574 => x"E3A02002",
000575 => x"E1A03002",
000576 => x"E5CD0010",
000577 => x"E1A01005",
000578 => x"E3A00072",
000579 => x"E58D4000",
000580 => x"EBFFFE6E",
000581 => x"E3A03002",
000582 => x"E5CD0011",
000583 => x"E1A01005",
000584 => x"E3A00072",
000585 => x"E3A02003",
000586 => x"E58D4000",
000587 => x"EBFFFE67",
000588 => x"E5DD300F",
000589 => x"E20000FF",
000590 => x"E3530053",
000591 => x"E5CD0012",
000592 => x"1A000002",
000593 => x"E5DD3010",
000594 => x"E353004D",
000595 => x"0A00006B",
000596 => x"E59F075C",
000597 => x"EBFFFEF4",
000598 => x"E3560000",
000599 => x"0AFFFFCD",
000600 => x"E59F0750",
000601 => x"EBFFFEF0",
000602 => x"E3A0100D",
000603 => x"E3A00000",
000604 => x"EBFFFED8",
000605 => x"E3A00006",
000606 => x"EBFFFEA0",
000607 => x"E3A01006",
000608 => x"E3C00008",
000609 => x"EBFFFED3",
000610 => x"E3A00006",
000611 => x"EBFFFE9B",
000612 => x"E1E00000",
000613 => x"E2000002",
000614 => x"E1E00000",
000615 => x"E3A01006",
000616 => x"EBFFFECC",
000617 => x"E3A00301",
000618 => x"EBFFFDAA",
000619 => x"EAFFFFFE",
000620 => x"E3540034",
000621 => x"0A000029",
000622 => x"CA00001C",
000623 => x"E3540031",
000624 => x"0A000036",
000625 => x"DA000098",
000626 => x"E3540032",
000627 => x"0A0000A2",
000628 => x"E3540033",
000629 => x"1A000098",
000630 => x"E1A00004",
000631 => x"EBFFFDFF",
000632 => x"E59F06D4",
000633 => x"EBFFFED0",
000634 => x"E1A00009",
000635 => x"E3A01002",
000636 => x"E3A02001",
000637 => x"EBFFFEDA",
000638 => x"E3A01002",
000639 => x"E1A00009",
000640 => x"EBFFFF3F",
000641 => x"E21010FF",
000642 => x"11A05001",
000643 => x"13A06000",
000644 => x"1AFFFFA8",
000645 => x"E59F06A4",
000646 => x"EBFFFEC3",
000647 => x"EAFFFF9D",
000648 => x"E3A04033",
000649 => x"E28DA006",
000650 => x"E28D900F",
000651 => x"EAFFFF9B",
000652 => x"E3540066",
000653 => x"0A00002A",
000654 => x"DA0000AD",
000655 => x"E3540068",
000656 => x"0A00010F",
000657 => x"E3540072",
000658 => x"1A00007B",
000659 => x"E1A00004",
000660 => x"EBFFFDE2",
000661 => x"E3A006FF",
000662 => x"E280F20F",
000663 => x"EAFFFFFE",
000664 => x"E1A00004",
000665 => x"EBFFFDDD",
000666 => x"E59F064C",
000667 => x"EBFFFEAE",
000668 => x"E1A00009",
000669 => x"E3A01002",
000670 => x"E3A02001",
000671 => x"EBFFFEB8",
000672 => x"E1A00009",
000673 => x"E3A01002",
000674 => x"EBFFFF1D",
000675 => x"E21080FF",
000676 => x"1A0000A4",
000677 => x"E59F0628",
000678 => x"EBFFFEA3",
000679 => x"EAFFFF7D",
000680 => x"E1A00004",
000681 => x"EBFFFDCD",
000682 => x"E59F0618",
000683 => x"EBFFFE9E",
000684 => x"E1A00009",
000685 => x"E3A01004",
000686 => x"E3A02000",
000687 => x"EBFFFEA8",
000688 => x"E5DD300F",
000689 => x"E3530053",
000690 => x"1A000002",
000691 => x"E5DD3010",
000692 => x"E353004D",
000693 => x"0A000115",
000694 => x"E59F05EC",
000695 => x"EBFFFE92",
000696 => x"EAFFFF6C",
000697 => x"E1A00004",
000698 => x"EBFFFDBC",
000699 => x"E59F05DC",
000700 => x"EBFFFE8D",
000701 => x"E59F05D8",
000702 => x"EBFFFE8B",
000703 => x"EAFFFF65",
000704 => x"E5DD3011",
000705 => x"E3530042",
000706 => x"1AFFFF90",
000707 => x"E3500052",
000708 => x"1AFFFF8E",
000709 => x"E1A01005",
000710 => x"E3A02004",
000711 => x"E2433040",
000712 => x"E2800020",
000713 => x"E58D4000",
000714 => x"EBFFFDE8",
000715 => x"E1A01005",
000716 => x"E5CD000F",
000717 => x"E3A02005",
000718 => x"E3A03002",
000719 => x"E3A00072",
000720 => x"E58D4000",
000721 => x"EBFFFDE1",
000722 => x"E1A01005",
000723 => x"E5CD0010",
000724 => x"E3A02006",
000725 => x"E3A03002",
000726 => x"E3A00072",
000727 => x"E58D4000",
000728 => x"EBFFFDDA",
000729 => x"E1A01005",
000730 => x"E5CD0011",
000731 => x"E3A02007",
000732 => x"E3A03002",
000733 => x"E3A00072",
000734 => x"E58D4000",
000735 => x"EBFFFDD3",
000736 => x"E5CD0012",
000737 => x"E1A00009",
000738 => x"EBFFFEF8",
000739 => x"E2907004",
000740 => x"0A000022",
000741 => x"E1A06004",
000742 => x"E2842008",
000743 => x"E1A01005",
000744 => x"E3A03002",
000745 => x"E3A00072",
000746 => x"E58D6000",
000747 => x"EBFFFDC7",
000748 => x"E2842009",
000749 => x"E5CD000F",
000750 => x"E1A01005",
000751 => x"E3A03002",
000752 => x"E3A00072",
000753 => x"E58D6000",
000754 => x"EBFFFDC0",
000755 => x"E284200A",
000756 => x"E5CD0010",
000757 => x"E1A01005",
000758 => x"E3A03002",
000759 => x"E3A00072",
000760 => x"E58D6000",
000761 => x"EBFFFDB9",
000762 => x"E284200B",
000763 => x"E5CD0011",
000764 => x"E1A01005",
000765 => x"E3A03002",
000766 => x"E3A00072",
000767 => x"E58D6000",
000768 => x"EBFFFDB2",
000769 => x"E5CD0012",
000770 => x"E1A00009",
000771 => x"EBFFFED7",
000772 => x"E4840004",
000773 => x"E1540007",
000774 => x"13540902",
000775 => x"3AFFFFDD",
000776 => x"E59F04B0",
000777 => x"EBFFFE40",
000778 => x"EAFFFF4C",
000779 => x"E3740001",
000780 => x"0AFFFF18",
000781 => x"E3540030",
000782 => x"0A000004",
000783 => x"E20400FF",
000784 => x"EBFFFD66",
000785 => x"E59F0490",
000786 => x"EBFFFE37",
000787 => x"EAFFFF11",
000788 => x"E1A00004",
000789 => x"EBFFFD61",
000790 => x"EAFFFF40",
000791 => x"E1A00004",
000792 => x"EBFFFD5E",
000793 => x"E59F0474",
000794 => x"EBFFFE2F",
000795 => x"EBFFFD55",
000796 => x"E3700001",
000797 => x"0AFFFFFC",
000798 => x"EBFFFD52",
000799 => x"E3700001",
000800 => x"1AFFFFFC",
000801 => x"E3A05301",
000802 => x"E5950000",
000803 => x"E1A0100A",
000804 => x"E3A02008",
000805 => x"EBFFFE52",
000806 => x"E5DD0006",
000807 => x"E3500000",
000808 => x"0A000005",
000809 => x"E3A04000",
000810 => x"E2844001",
000811 => x"EBFFFD4B",
000812 => x"E7D4000A",
000813 => x"E3500000",
000814 => x"1AFFFFFA",
000815 => x"E3A00020",
000816 => x"EBFFFD46",
000817 => x"EBFFFD3F",
000818 => x"E3700001",
000819 => x"1A000005",
000820 => x"E3A03301",
000821 => x"E2833E9E",
000822 => x"E2855004",
000823 => x"E2833004",
000824 => x"E1550003",
000825 => x"1AFFFFE7",
000826 => x"E59F03F4",
000827 => x"EBFFFE0E",
000828 => x"EAFFFEE8",
000829 => x"E3540035",
000830 => x"0A0000AE",
000831 => x"E3540061",
000832 => x"1AFFFFCD",
000833 => x"E1A00004",
000834 => x"EBFFFD34",
000835 => x"E59F03D4",
000836 => x"EBFFFE05",
000837 => x"E59F03D0",
000838 => x"EBFFFE03",
000839 => x"E59F03CC",
000840 => x"EBFFFE01",
000841 => x"EAFFFEDB",
000842 => x"E59F03C4",
000843 => x"EBFFFDFE",
000844 => x"E1A00009",
000845 => x"E3A01004",
000846 => x"E3A02000",
000847 => x"EBFFFE08",
000848 => x"E5DD300F",
000849 => x"E3530053",
000850 => x"1A000002",
000851 => x"E5DD2010",
000852 => x"E352004D",
000853 => x"0A000004",
000854 => x"E59F0398",
000855 => x"EBFFFDF2",
000856 => x"E59F0394",
000857 => x"EBFFFDF0",
000858 => x"EAFFFECA",
000859 => x"E5DD1011",
000860 => x"E3510042",
000861 => x"1AFFFFF7",
000862 => x"E5DD0012",
000863 => x"E3500052",
000864 => x"1AFFFFF4",
000865 => x"E3A04000",
000866 => x"E5C43000",
000867 => x"E1A00000",
000868 => x"E5C42001",
000869 => x"E1A00000",
000870 => x"E5C41002",
000871 => x"E1A00000",
000872 => x"E5C40003",
000873 => x"E1A00000",
000874 => x"E241103E",
000875 => x"E1A00009",
000876 => x"E1A02004",
000877 => x"EBFFFDEA",
000878 => x"E5DD300F",
000879 => x"E5C43004",
000880 => x"E5DD2010",
000881 => x"E5C42005",
000882 => x"E5DD3011",
000883 => x"E5C43006",
000884 => x"E5DD2012",
000885 => x"E1A00009",
000886 => x"E5C42007",
000887 => x"EBFFFE63",
000888 => x"E3A03CFF",
000889 => x"E28330FC",
000890 => x"E1500003",
000891 => x"E1A05000",
000892 => x"8A00009A",
000893 => x"E3700004",
000894 => x"12844008",
000895 => x"1280600B",
000896 => x"0A000006",
000897 => x"EBFFFCEF",
000898 => x"E3700001",
000899 => x"0AFFFFFC",
000900 => x"E1560004",
000901 => x"E5C40000",
000902 => x"E2844001",
000903 => x"1AFFFFF8",
000904 => x"E59F02D8",
000905 => x"EBFFFDC0",
000906 => x"E59F02D4",
000907 => x"EBFFFDBE",
000908 => x"E375000C",
000909 => x"0A00000F",
000910 => x"E3A04000",
000911 => x"E285700C",
000912 => x"E1A06004",
000913 => x"E5D45000",
000914 => x"E3A00077",
000915 => x"E1A01008",
000916 => x"E1A02006",
000917 => x"E3A03002",
000918 => x"E58D5000",
000919 => x"EBFFFD1B",
000920 => x"E3500000",
000921 => x"1AFFFFF7",
000922 => x"E2844001",
000923 => x"E1540007",
000924 => x"E1A06004",
000925 => x"1AFFFFF2",
000926 => x"E59F0288",
000927 => x"EBFFFDAA",
000928 => x"EAFFFFB6",
000929 => x"E1A00004",
000930 => x"EBFFFCD4",
000931 => x"E59F0278",
000932 => x"EBFFFDA5",
000933 => x"E59F0274",
000934 => x"EBFFFDA3",
000935 => x"E59F0270",
000936 => x"EBFFFDA1",
000937 => x"E59F026C",
000938 => x"EBFFFD9F",
000939 => x"E59F0268",
000940 => x"EBFFFD9D",
000941 => x"E59F0264",
000942 => x"EBFFFD9B",
000943 => x"E59F0260",
000944 => x"EBFFFD99",
000945 => x"E59F025C",
000946 => x"EBFFFD97",
000947 => x"E59F0258",
000948 => x"EBFFFD95",
000949 => x"E59F0254",
000950 => x"EBFFFD93",
000951 => x"E59F0250",
000952 => x"EBFFFD91",
000953 => x"E59F024C",
000954 => x"EBFFFD8F",
000955 => x"E59F0248",
000956 => x"EBFFFD8D",
000957 => x"E59F0244",
000958 => x"EBFFFD8B",
000959 => x"E59F0240",
000960 => x"EBFFFD89",
000961 => x"E59F023C",
000962 => x"EBFFFD87",
000963 => x"E59F0238",
000964 => x"EBFFFD85",
000965 => x"E59F0234",
000966 => x"EBFFFD83",
000967 => x"E59F0230",
000968 => x"EBFFFD81",
000969 => x"E59F022C",
000970 => x"EBFFFD7F",
000971 => x"EAFFFE59",
000972 => x"E5DD3011",
000973 => x"E3530042",
000974 => x"1AFFFEE6",
000975 => x"E5DD3012",
000976 => x"E3530052",
000977 => x"1AFFFEE3",
000978 => x"E3A01004",
000979 => x"E3A02000",
000980 => x"E1A00009",
000981 => x"EBFFFD82",
000982 => x"E1A00009",
000983 => x"EBFFFE03",
000984 => x"E3A03C7F",
000985 => x"E28330F8",
000986 => x"E1500003",
000987 => x"8A00003B",
000988 => x"E2804301",
000989 => x"E2844004",
000990 => x"E3540301",
000991 => x"0A000009",
000992 => x"E3A05301",
000993 => x"E3A01004",
000994 => x"E3A02000",
000995 => x"E1A00009",
000996 => x"EBFFFD73",
000997 => x"E1A00009",
000998 => x"EBFFFDF4",
000999 => x"E4850004",
001000 => x"E1550004",
001001 => x"1AFFFFF6",
001002 => x"E59F00FC",
001003 => x"EBFFFD5E",
001004 => x"EBFFFDF6",
001005 => x"EAFFFE37",
001006 => x"E1A00004",
001007 => x"EBFFFC87",
001008 => x"E59F0194",
001009 => x"EBFFFD58",
001010 => x"E1A00009",
001011 => x"E3A01002",
001012 => x"E3A02001",
001013 => x"EBFFFD62",
001014 => x"E1A00009",
001015 => x"E3A01002",
001016 => x"EBFFFDC7",
001017 => x"E21060FF",
001018 => x"0AFFFE89",
001019 => x"E59F016C",
001020 => x"EBFFFD4D",
001021 => x"E59F0168",
001022 => x"EBFFFD4B",
001023 => x"EBFFFC71",
001024 => x"E3700001",
001025 => x"0AFFFFFC",
001026 => x"EBFFFC6E",
001027 => x"E3700001",
001028 => x"1AFFFFFC",
001029 => x"E3A05000",
001030 => x"EA000001",
001031 => x"E3540000",
001032 => x"AA000011",
001033 => x"E3A0C000",
001034 => x"E1A02005",
001035 => x"E1A01006",
001036 => x"E3A03002",
001037 => x"E3A00072",
001038 => x"E58DC000",
001039 => x"EBFFFCA3",
001040 => x"E1A04000",
001041 => x"EBFFFC5F",
001042 => x"E3700001",
001043 => x"E1A00004",
001044 => x"0AFFFFF1",
001045 => x"E59F010C",
001046 => x"EBFFFD33",
001047 => x"EAFFFF21",
001048 => x"E59F0104",
001049 => x"EBFFFD30",
001050 => x"EAFFFE0A",
001051 => x"EBFFFC5B",
001052 => x"E3A03801",
001053 => x"E2855001",
001054 => x"E2433001",
001055 => x"E1550003",
001056 => x"1AFFFFE7",
001057 => x"EAFFFF17",
001058 => x"000112AC",
001059 => x"000112F8",
001060 => x"00011340",
001061 => x"00011388",
001062 => x"000113D0",
001063 => x"00011418",
001064 => x"00011460",
001065 => x"000114CC",
001066 => x"00011504",
001067 => x"00011514",
001068 => x"000116A0",
001069 => x"00011704",
001070 => x"00011E08",
001071 => x"00011644",
001072 => x"00011680",
001073 => x"00011730",
001074 => x"00011518",
001075 => x"000115B0",
001076 => x"00011D8C",
001077 => x"00011DBC",
001078 => x"000116F0",
001079 => x"00011DE4",
001080 => x"000115D8",
001081 => x"00011620",
001082 => x"000118E0",
001083 => x"00011914",
001084 => x"00011980",
001085 => x"00011750",
001086 => x"000117F8",
001087 => x"00011DD8",
001088 => x"000117B0",
001089 => x"000117C8",
001090 => x"000117E8",
001091 => x"000119C4",
001092 => x"000119E0",
001093 => x"00011A00",
001094 => x"00011A40",
001095 => x"00011A74",
001096 => x"00011AB0",
001097 => x"00011AEC",
001098 => x"00011B10",
001099 => x"00011B4C",
001100 => x"00011B68",
001101 => x"00011B80",
001102 => x"00011BC8",
001103 => x"00011C08",
001104 => x"00011C40",
001105 => x"00011C64",
001106 => x"00011CA8",
001107 => x"00011CE8",
001108 => x"00011D14",
001109 => x"00011D40",
001110 => x"00011D64",
001111 => x"0001181C",
001112 => x"00011858",
001113 => x"00011898",
001114 => x"00011E2C",
001115 => x"0001158C",
001116 => x"E10F3000",
001117 => x"E3C330C0",
001118 => x"E129F003",
001119 => x"E1A0F00E",
001120 => x"E10F3000",
001121 => x"E38330C0",
001122 => x"E129F003",
001123 => x"E1A0F00E",
001124 => x"00000000",
001125 => x"2030202D",
001126 => x"20626F6F",
001127 => x"74206672",
001128 => x"6F6D2063",
001129 => x"6F726520",
001130 => x"52414D20",
001131 => x"28737461",
001132 => x"72742061",
001133 => x"70706C69",
001134 => x"63617469",
001135 => x"6F6E290D",
001136 => x"0A203120",
001137 => x"2D207072",
001138 => x"6F677261",
001139 => x"6D20636F",
001140 => x"72652052",
001141 => x"414D2076",
001142 => x"69612055",
001143 => x"4152545F",
001144 => x"300D0A20",
001145 => x"32202D20",
001146 => x"636F7265",
001147 => x"2052414D",
001148 => x"2064756D",
001149 => x"700D0A00",
001150 => x"2033202D",
001151 => x"20626F6F",
001152 => x"74206672",
001153 => x"6F6D2049",
001154 => x"32432045",
001155 => x"4550524F",
001156 => x"4D0D0A20",
001157 => x"34202D20",
001158 => x"70726F67",
001159 => x"72616D20",
001160 => x"49324320",
001161 => x"45455052",
001162 => x"4F4D2076",
001163 => x"69612055",
001164 => x"4152545F",
001165 => x"300D0A20",
001166 => x"35202D20",
001167 => x"73686F77",
001168 => x"20636F6E",
001169 => x"74656E74",
001170 => x"206F6620",
001171 => x"49324320",
001172 => x"45455052",
001173 => x"4F4D0D0A",
001174 => x"00000000",
001175 => x"2061202D",
001176 => x"20617574",
001177 => x"6F6D6174",
001178 => x"69632062",
001179 => x"6F6F7420",
001180 => x"636F6E66",
001181 => x"69677572",
001182 => x"6174696F",
001183 => x"6E0D0A20",
001184 => x"68202D20",
001185 => x"68656C70",
001186 => x"0D0A2072",
001187 => x"202D2072",
001188 => x"65737461",
001189 => x"72742073",
001190 => x"79737465",
001191 => x"6D0D0A0D",
001192 => x"0A53656C",
001193 => x"6563743A",
001194 => x"20000000",
001195 => x"0D0A0D0A",
001196 => x"0D0A2B2D",
001197 => x"2D2D2D2D",
001198 => x"2D2D2D2D",
001199 => x"2D2D2D2D",
001200 => x"2D2D2D2D",
001201 => x"2D2D2D2D",
001202 => x"2D2D2D2D",
001203 => x"2D2D2D2D",
001204 => x"2D2D2D2D",
001205 => x"2D2D2D2D",
001206 => x"2D2D2D2D",
001207 => x"2D2D2D2D",
001208 => x"2D2D2D2D",
001209 => x"2D2D2D2D",
001210 => x"2D2D2D2D",
001211 => x"2D2D2D2D",
001212 => x"2D2D2D2B",
001213 => x"0D0A0000",
001214 => x"7C202020",
001215 => x"203C3C3C",
001216 => x"2053544F",
001217 => x"524D2043",
001218 => x"6F726520",
001219 => x"50726F63",
001220 => x"6573736F",
001221 => x"72205379",
001222 => x"7374656D",
001223 => x"202D2042",
001224 => x"79205374",
001225 => x"65706861",
001226 => x"6E204E6F",
001227 => x"6C74696E",
001228 => x"67203E3E",
001229 => x"3E202020",
001230 => x"207C0D0A",
001231 => x"00000000",
001232 => x"2B2D2D2D",
001233 => x"2D2D2D2D",
001234 => x"2D2D2D2D",
001235 => x"2D2D2D2D",
001236 => x"2D2D2D2D",
001237 => x"2D2D2D2D",
001238 => x"2D2D2D2D",
001239 => x"2D2D2D2D",
001240 => x"2D2D2D2D",
001241 => x"2D2D2D2D",
001242 => x"2D2D2D2D",
001243 => x"2D2D2D2D",
001244 => x"2D2D2D2D",
001245 => x"2D2D2D2D",
001246 => x"2D2D2D2D",
001247 => x"2D2D2D2D",
001248 => x"2D2B0D0A",
001249 => x"00000000",
001250 => x"7C202020",
001251 => x"20202020",
001252 => x"2020426F",
001253 => x"6F746C6F",
001254 => x"61646572",
001255 => x"20666F72",
001256 => x"2053544F",
001257 => x"524D2053",
001258 => x"6F432020",
001259 => x"20566572",
001260 => x"73696F6E",
001261 => x"3A203230",
001262 => x"31323035",
001263 => x"32342D44",
001264 => x"20202020",
001265 => x"20202020",
001266 => x"207C0D0A",
001267 => x"00000000",
001268 => x"7C202020",
001269 => x"20202020",
001270 => x"20202020",
001271 => x"20202020",
001272 => x"436F6E74",
001273 => x"6163743A",
001274 => x"2073746E",
001275 => x"6F6C7469",
001276 => x"6E674067",
001277 => x"6F6F676C",
001278 => x"656D6169",
001279 => x"6C2E636F",
001280 => x"6D202020",
001281 => x"20202020",
001282 => x"20202020",
001283 => x"20202020",
001284 => x"207C0D0A",
001285 => x"00000000",
001286 => x"2B2D2D2D",
001287 => x"2D2D2D2D",
001288 => x"2D2D2D2D",
001289 => x"2D2D2D2D",
001290 => x"2D2D2D2D",
001291 => x"2D2D2D2D",
001292 => x"2D2D2D2D",
001293 => x"2D2D2D2D",
001294 => x"2D2D2D2D",
001295 => x"2D2D2D2D",
001296 => x"2D2D2D2D",
001297 => x"2D2D2D2D",
001298 => x"2D2D2D2D",
001299 => x"2D2D2D2D",
001300 => x"2D2D2D2D",
001301 => x"2D2D2D2D",
001302 => x"2D2B0D0A",
001303 => x"0D0A0000",
001304 => x"203C2057",
001305 => x"656C636F",
001306 => x"6D652074",
001307 => x"6F207468",
001308 => x"65205354",
001309 => x"4F524D20",
001310 => x"536F4320",
001311 => x"626F6F74",
001312 => x"6C6F6164",
001313 => x"65722063",
001314 => x"6F6E736F",
001315 => x"6C652120",
001316 => x"3E0D0A20",
001317 => x"3C205365",
001318 => x"6C656374",
001319 => x"20616E20",
001320 => x"6F706572",
001321 => x"6174696F",
001322 => x"6E206672",
001323 => x"6F6D2074",
001324 => x"6865206D",
001325 => x"656E7520",
001326 => x"62656C6F",
001327 => x"77206F72",
001328 => x"20707265",
001329 => x"7373203E",
001330 => x"0D0A0000",
001331 => x"203C2074",
001332 => x"68652062",
001333 => x"6F6F7420",
001334 => x"6B657920",
001335 => x"666F7220",
001336 => x"696D6D65",
001337 => x"64696174",
001338 => x"65206170",
001339 => x"706C6963",
001340 => x"6174696F",
001341 => x"6E207374",
001342 => x"6172742E",
001343 => x"203E0D0A",
001344 => x"0D0A0000",
001345 => x"204C6F61",
001346 => x"64204164",
001347 => x"64726573",
001348 => x"733A2000",
001349 => x"0A0D0000",
001350 => x"0D0A0D0A",
001351 => x"4170706C",
001352 => x"69636174",
001353 => x"696F6E20",
001354 => x"77696C6C",
001355 => x"20737461",
001356 => x"72742061",
001357 => x"75746F6D",
001358 => x"61746963",
001359 => x"616C6C79",
001360 => x"20616674",
001361 => x"65722064",
001362 => x"6F776E6C",
001363 => x"6F61642E",
001364 => x"0D0A2D3E",
001365 => x"20576169",
001366 => x"74696E67",
001367 => x"20666F72",
001368 => x"20277374",
001369 => x"6F726D5F",
001370 => x"70726F67",
001371 => x"72616D2E",
001372 => x"62696E27",
001373 => x"20696E20",
001374 => x"62797465",
001375 => x"2D737472",
001376 => x"65616D20",
001377 => x"6D6F6465",
001378 => x"2E2E2E00",
001379 => x"20455252",
001380 => x"4F522120",
001381 => x"50726F67",
001382 => x"72616D20",
001383 => x"66696C65",
001384 => x"20746F6F",
001385 => x"20626967",
001386 => x"210D0A0D",
001387 => x"0A000000",
001388 => x"20496E76",
001389 => x"616C6964",
001390 => x"2070726F",
001391 => x"6772616D",
001392 => x"6D696E67",
001393 => x"2066696C",
001394 => x"65210D0A",
001395 => x"0D0A5365",
001396 => x"6C656374",
001397 => x"3A200000",
001398 => x"0D0A0D0A",
001399 => x"41626F72",
001400 => x"74206475",
001401 => x"6D70696E",
001402 => x"67206279",
001403 => x"20707265",
001404 => x"7373696E",
001405 => x"6720616E",
001406 => x"79206B65",
001407 => x"792E0D0A",
001408 => x"50726573",
001409 => x"7320616E",
001410 => x"79206B65",
001411 => x"7920746F",
001412 => x"20636F6E",
001413 => x"74696E75",
001414 => x"652E0D0A",
001415 => x"0D0A0000",
001416 => x"0D0A0D0A",
001417 => x"44756D70",
001418 => x"696E6720",
001419 => x"636F6D70",
001420 => x"6C657465",
001421 => x"642E0D0A",
001422 => x"0D0A5365",
001423 => x"6C656374",
001424 => x"3A200000",
001425 => x"0D0A0D0A",
001426 => x"456E7465",
001427 => x"72206465",
001428 => x"76696365",
001429 => x"20616464",
001430 => x"72657373",
001431 => x"20283278",
001432 => x"20686578",
001433 => x"5F636861",
001434 => x"72732C20",
001435 => x"73657420",
001436 => x"4C534220",
001437 => x"746F2027",
001438 => x"3027293A",
001439 => x"20000000",
001440 => x"20496E76",
001441 => x"616C6964",
001442 => x"20616464",
001443 => x"72657373",
001444 => x"210D0A0D",
001445 => x"0A53656C",
001446 => x"6563743A",
001447 => x"20000000",
001448 => x"0D0A4170",
001449 => x"706C6963",
001450 => x"6174696F",
001451 => x"6E207769",
001452 => x"6C6C2073",
001453 => x"74617274",
001454 => x"20617574",
001455 => x"6F6D6174",
001456 => x"6963616C",
001457 => x"6C792061",
001458 => x"66746572",
001459 => x"2075706C",
001460 => x"6F61642E",
001461 => x"0D0A2D3E",
001462 => x"204C6F61",
001463 => x"64696E67",
001464 => x"20626F6F",
001465 => x"7420696D",
001466 => x"6167652E",
001467 => x"2E2E0000",
001468 => x"2055706C",
001469 => x"6F616420",
001470 => x"636F6D70",
001471 => x"6C657465",
001472 => x"0D0A0000",
001473 => x"20496E76",
001474 => x"616C6964",
001475 => x"20626F6F",
001476 => x"74206465",
001477 => x"76696365",
001478 => x"206F7220",
001479 => x"66696C65",
001480 => x"210D0A0D",
001481 => x"0A53656C",
001482 => x"6563743A",
001483 => x"20000000",
001484 => x"0D0A496E",
001485 => x"76616C69",
001486 => x"64206164",
001487 => x"64726573",
001488 => x"73210D0A",
001489 => x"0D0A5365",
001490 => x"6C656374",
001491 => x"3A200000",
001492 => x"0D0A4461",
001493 => x"74612077",
001494 => x"696C6C20",
001495 => x"6F766572",
001496 => x"77726974",
001497 => x"65205241",
001498 => x"4D20636F",
001499 => x"6E74656E",
001500 => x"74210D0A",
001501 => x"2D3E2057",
001502 => x"61697469",
001503 => x"6E672066",
001504 => x"6F722027",
001505 => x"73746F72",
001506 => x"6D5F7072",
001507 => x"6F677261",
001508 => x"6D2E6269",
001509 => x"6E272069",
001510 => x"6E206279",
001511 => x"74652D73",
001512 => x"74726561",
001513 => x"6D206D6F",
001514 => x"64652E2E",
001515 => x"2E000000",
001516 => x"20446F77",
001517 => x"6E6C6F61",
001518 => x"6420636F",
001519 => x"6D706C65",
001520 => x"7465640D",
001521 => x"0A000000",
001522 => x"57726974",
001523 => x"696E6720",
001524 => x"62756666",
001525 => x"65722074",
001526 => x"6F206932",
001527 => x"63204545",
001528 => x"50524F4D",
001529 => x"2E2E2E00",
001530 => x"20436F6D",
001531 => x"706C6574",
001532 => x"65640D0A",
001533 => x"0D0A0000",
001534 => x"20496E76",
001535 => x"616C6964",
001536 => x"20626F6F",
001537 => x"74206465",
001538 => x"76696365",
001539 => x"206F7220",
001540 => x"66696C65",
001541 => x"210D0A0D",
001542 => x"0A000000",
001543 => x"0D0A0D0A",
001544 => x"456E7465",
001545 => x"72206465",
001546 => x"76696365",
001547 => x"20616464",
001548 => x"72657373",
001549 => x"20283220",
001550 => x"6865782D",
001551 => x"63686172",
001552 => x"732C2073",
001553 => x"6574204C",
001554 => x"53422074",
001555 => x"6F202730",
001556 => x"27293A20",
001557 => x"00000000",
001558 => x"0D0A0D0A",
001559 => x"41626F72",
001560 => x"74206475",
001561 => x"6D70696E",
001562 => x"67206279",
001563 => x"20707265",
001564 => x"7373696E",
001565 => x"6720616E",
001566 => x"79206B65",
001567 => x"792E2049",
001568 => x"66206E6F",
001569 => x"20646174",
001570 => x"61206973",
001571 => x"2073686F",
001572 => x"776E2C0D",
001573 => x"0A000000",
001574 => x"74686520",
001575 => x"73656C65",
001576 => x"63746564",
001577 => x"20646576",
001578 => x"69636520",
001579 => x"6973206E",
001580 => x"6F742072",
001581 => x"6573706F",
001582 => x"6E64696E",
001583 => x"672E2050",
001584 => x"72657373",
001585 => x"20616E79",
001586 => x"206B6579",
001587 => x"20746F20",
001588 => x"636F6E74",
001589 => x"696E7565",
001590 => x"2E0D0A0D",
001591 => x"0A000000",
001592 => x"0D0A0D0A",
001593 => x"4175746F",
001594 => x"6D617469",
001595 => x"6320626F",
001596 => x"6F742063",
001597 => x"6F6E6669",
001598 => x"67757261",
001599 => x"74696F6E",
001600 => x"20666F72",
001601 => x"20706F77",
001602 => x"65722D75",
001603 => x"703A0D0A",
001604 => x"00000000",
001605 => x"5B333231",
001606 => x"305D2063",
001607 => x"6F6E6669",
001608 => x"67757261",
001609 => x"74696F6E",
001610 => x"20444950",
001611 => x"20737769",
001612 => x"7463680D",
001613 => x"0A203030",
001614 => x"3030202D",
001615 => x"20537461",
001616 => x"72742062",
001617 => x"6F6F746C",
001618 => x"6F616465",
001619 => x"7220636F",
001620 => x"6E736F6C",
001621 => x"650D0A20",
001622 => x"30303031",
001623 => x"202D2041",
001624 => x"75746F6D",
001625 => x"61746963",
001626 => x"20626F6F",
001627 => x"74206672",
001628 => x"6F6D2063",
001629 => x"6F726520",
001630 => x"52414D0D",
001631 => x"0A000000",
001632 => x"20303031",
001633 => x"30202D20",
001634 => x"4175746F",
001635 => x"6D617469",
001636 => x"6320626F",
001637 => x"6F742066",
001638 => x"726F6D20",
001639 => x"49324320",
001640 => x"45455052",
001641 => x"4F4D2028",
001642 => x"41646472",
001643 => x"65737320",
001644 => x"30784130",
001645 => x"290D0A0D",
001646 => x"0A53656C",
001647 => x"6563743A",
001648 => x"20000000",
001649 => x"0D0A0D0A",
001650 => x"53544F52",
001651 => x"4D20536F",
001652 => x"4320626F",
001653 => x"6F746C6F",
001654 => x"61646572",
001655 => x"0D0A0000",
001656 => x"2730273A",
001657 => x"20457865",
001658 => x"63757465",
001659 => x"2070726F",
001660 => x"6772616D",
001661 => x"20696E20",
001662 => x"52414D2E",
001663 => x"0D0A0000",
001664 => x"2731273A",
001665 => x"20577269",
001666 => x"74652027",
001667 => x"73746F72",
001668 => x"6D5F7072",
001669 => x"6F677261",
001670 => x"6D2E6269",
001671 => x"6E272074",
001672 => x"6F207468",
001673 => x"6520636F",
001674 => x"72652773",
001675 => x"2052414D",
001676 => x"20766961",
001677 => x"20554152",
001678 => x"542E0D0A",
001679 => x"00000000",
001680 => x"2732273A",
001681 => x"20507269",
001682 => x"6E742063",
001683 => x"75727265",
001684 => x"6E742063",
001685 => x"6F6E7465",
001686 => x"6E74206F",
001687 => x"6620636F",
001688 => x"6D706C65",
001689 => x"74652063",
001690 => x"6F726520",
001691 => x"52414D2E",
001692 => x"0D0A0000",
001693 => x"2733273A",
001694 => x"204C6F61",
001695 => x"6420626F",
001696 => x"6F742069",
001697 => x"6D616765",
001698 => x"2066726F",
001699 => x"6D204545",
001700 => x"50524F4D",
001701 => x"20616E64",
001702 => x"20737461",
001703 => x"72742061",
001704 => x"70706C69",
001705 => x"63617469",
001706 => x"6F6E2E0D",
001707 => x"0A000000",
001708 => x"2734273A",
001709 => x"20577269",
001710 => x"74652027",
001711 => x"73746F72",
001712 => x"6D5F7072",
001713 => x"6F677261",
001714 => x"6D2E6269",
001715 => x"6E272074",
001716 => x"6F204932",
001717 => x"43204545",
001718 => x"50524F4D",
001719 => x"20766961",
001720 => x"20554152",
001721 => x"542E0D0A",
001722 => x"00000000",
001723 => x"2735273A",
001724 => x"20507269",
001725 => x"6E742063",
001726 => x"6F6E7465",
001727 => x"6E74206F",
001728 => x"66204932",
001729 => x"43204545",
001730 => x"50524F4D",
001731 => x"2E0D0A00",
001732 => x"2761273A",
001733 => x"2053686F",
001734 => x"77204449",
001735 => x"50207377",
001736 => x"69746368",
001737 => x"20636F6E",
001738 => x"66696775",
001739 => x"72617469",
001740 => x"6F6E7320",
001741 => x"666F7220",
001742 => x"6175746F",
001743 => x"6D617469",
001744 => x"6320626F",
001745 => x"6F742E0D",
001746 => x"0A000000",
001747 => x"2768273A",
001748 => x"2053686F",
001749 => x"77207468",
001750 => x"69732073",
001751 => x"63726565",
001752 => x"6E2E0D0A",
001753 => x"00000000",
001754 => x"2772273A",
001755 => x"20526573",
001756 => x"65742073",
001757 => x"79737465",
001758 => x"6D2E0D0A",
001759 => x"0D0A0000",
001760 => x"426F6F74",
001761 => x"20454550",
001762 => x"524F4D3A",
001763 => x"20323478",
001764 => x"786E6E6E",
001765 => x"20286C69",
001766 => x"6B652032",
001767 => x"34414136",
001768 => x"34292C20",
001769 => x"37206269",
001770 => x"74206164",
001771 => x"64726573",
001772 => x"73202B20",
001773 => x"646F6E74",
001774 => x"2D636172",
001775 => x"65206269",
001776 => x"742C0D0A",
001777 => x"00000000",
001778 => x"636F6E6E",
001779 => x"65637465",
001780 => x"6420746F",
001781 => x"20493243",
001782 => x"5F434F4E",
001783 => x"54524F4C",
001784 => x"4C45525F",
001785 => x"302C206F",
001786 => x"70657261",
001787 => x"74696E67",
001788 => x"20667265",
001789 => x"7175656E",
001790 => x"63792069",
001791 => x"73203130",
001792 => x"306B487A",
001793 => x"2C0D0A00",
001794 => x"6D617869",
001795 => x"6D756D20",
001796 => x"45455052",
001797 => x"4F4D2073",
001798 => x"697A6520",
001799 => x"3D203635",
001800 => x"35333620",
001801 => x"62797465",
001802 => x"203D3E20",
001803 => x"31362062",
001804 => x"69742061",
001805 => x"64647265",
001806 => x"73736573",
001807 => x"2C0D0A00",
001808 => x"66697865",
001809 => x"6420626F",
001810 => x"6F742064",
001811 => x"65766963",
001812 => x"65206164",
001813 => x"64726573",
001814 => x"733A2030",
001815 => x"7841300D",
001816 => x"0A0D0A00",
001817 => x"5465726D",
001818 => x"696E616C",
001819 => x"20736574",
001820 => x"75703A20",
001821 => x"39363030",
001822 => x"20626175",
001823 => x"642C2038",
001824 => x"20646174",
001825 => x"61206269",
001826 => x"74732C20",
001827 => x"6E6F2070",
001828 => x"61726974",
001829 => x"792C2031",
001830 => x"2073746F",
001831 => x"70206269",
001832 => x"740D0A0D",
001833 => x"0A000000",
001834 => x"466F7220",
001835 => x"6D6F7265",
001836 => x"20696E66",
001837 => x"6F726D61",
001838 => x"74696F6E",
001839 => x"20736565",
001840 => x"20746865",
001841 => x"2053544F",
001842 => x"524D2043",
001843 => x"6F726520",
001844 => x"2F205354",
001845 => x"4F524D20",
001846 => x"536F4320",
001847 => x"64617461",
001848 => x"73686565",
001849 => x"740D0A00",
001850 => x"68747470",
001851 => x"3A2F2F6F",
001852 => x"70656E63",
001853 => x"6F726573",
001854 => x"2E6F7267",
001855 => x"2F70726F",
001856 => x"6A656374",
001857 => x"2C73746F",
001858 => x"726D5F63",
001859 => x"6F72650D",
001860 => x"0A000000",
001861 => x"68747470",
001862 => x"3A2F2F6F",
001863 => x"70656E63",
001864 => x"6F726573",
001865 => x"2E6F7267",
001866 => x"2F70726F",
001867 => x"6A656374",
001868 => x"2C73746F",
001869 => x"726D5F73",
001870 => x"6F630D0A",
001871 => x"00000000",
001872 => x"436F6E74",
001873 => x"6163743A",
001874 => x"2073746E",
001875 => x"6F6C7469",
001876 => x"6E674067",
001877 => x"6F6F676C",
001878 => x"656D6169",
001879 => x"6C2E636F",
001880 => x"6D0D0A00",
001881 => x"28632920",
001882 => x"32303132",
001883 => x"20627920",
001884 => x"53746570",
001885 => x"68616E20",
001886 => x"4E6F6C74",
001887 => x"696E670D",
001888 => x"0A0D0A53",
001889 => x"656C6563",
001890 => x"743A2000",
001891 => x"0D0A0D0A",
001892 => x"5765276C",
001893 => x"6C207365",
001894 => x"6E642079",
001895 => x"6F752062",
001896 => x"61636B20",
001897 => x"2D20746F",
001898 => x"20746865",
001899 => x"20667574",
001900 => x"75726521",
001901 => x"2E0D0A0D",
001902 => x"0A000000",
001903 => x"202D2044",
001904 => x"6F63746F",
001905 => x"7220456D",
001906 => x"6D657420",
001907 => x"4C2E2042",
001908 => x"726F776E",
001909 => x"0D0A0D0A",
001910 => x"53656C65",
001911 => x"63743A20",
001912 => x"00000000",
001913 => x"20496E76",
001914 => x"616C6964",
001915 => x"206F7065",
001916 => x"72617469",
001917 => x"6F6E210D",
001918 => x"0A547279",
001919 => x"20616761",
001920 => x"696E3A20",
001921 => x"00000000",
001922 => x"0D0A0D0A",
001923 => x"2D3E2053",
001924 => x"74617274",
001925 => x"696E6720",
001926 => x"6170706C",
001927 => x"69636174",
001928 => x"696F6E2E",
001929 => x"2E2E0D0A",
001930 => x"0D0A0000",
001931 => x"0D0A0D0A",
001932 => x"41626F72",
001933 => x"74656421",
001934 => x"00000000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;