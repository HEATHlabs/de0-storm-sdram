-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
--				MEM_SIZE      : natural := 1024;  -- memory cells
--				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				MEM_SIZE      : natural := 2048;  -- memory cells
				LOG2_MEM_SIZE : natural := 11;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
	--bootloader_sdram
000000 => x"EA000006",
000001 => x"EAFFFFFE",
000002 => x"EAFFFFFE",
000003 => x"EAFFFFFE",
000004 => x"EAFFFFFE",
000005 => x"E1A00000",
000006 => x"EAFFFFFE",
000007 => x"EAFFFFFE",
000008 => x"E59F0034",
000009 => x"E10F1000",
000010 => x"E3C1107F",
000011 => x"E38110DF",
000012 => x"E129F001",
000013 => x"E1A0D000",
000014 => x"E3A00000",
000015 => x"E1A01000",
000016 => x"E1A02000",
000017 => x"E1A0B000",
000018 => x"E1A07000",
000019 => x"E59FA00C",
000020 => x"E1A0E00F",
000021 => x"E1A0F00A",
000022 => x"EAFFFFFE",
000023 => x"00002000",
000024 => x"00010784",
000025 => x"E3E03A0F",
000026 => x"E5131FFB",
000027 => x"E20020FF",
000028 => x"E3A00001",
000029 => x"E0010210",
000030 => x"E1A0F00E",
000031 => x"E3E03A0F",
000032 => x"E5130FFB",
000033 => x"E1A0F00E",
000034 => x"E3E01A0F",
000035 => x"E5113FFF",
000036 => x"E20000FF",
000037 => x"E3A02001",
000038 => x"E1833012",
000039 => x"E5013FFF",
000040 => x"E1A0F00E",
000041 => x"E20000FF",
000042 => x"E3A02001",
000043 => x"E1A02012",
000044 => x"E3E01A0F",
000045 => x"E5113FFF",
000046 => x"E1E02002",
000047 => x"E0033002",
000048 => x"E5013FFF",
000049 => x"E1A0F00E",
000050 => x"E3E01A0F",
000051 => x"E5113FFF",
000052 => x"E20000FF",
000053 => x"E3A02001",
000054 => x"E0233012",
000055 => x"E5013FFF",
000056 => x"E1A0F00E",
000057 => x"E3E03A0F",
000058 => x"E5030FFF",
000059 => x"E1A0F00E",
000060 => x"E20000FF",
000061 => x"E3500007",
000062 => x"E92D4010",
000063 => x"E3A0C000",
000064 => x"E3E0E0FF",
000065 => x"E20110FF",
000066 => x"8A000011",
000067 => x"E2403004",
000068 => x"E20330FF",
000069 => x"E3500003",
000070 => x"E1A0E183",
000071 => x"E3E04A0F",
000072 => x"E1A0C180",
000073 => x"9A000007",
000074 => x"E3A030FF",
000075 => x"E1A03E13",
000076 => x"E5142F8B",
000077 => x"E1E03003",
000078 => x"E0022003",
000079 => x"E1822E11",
000080 => x"E5042F8B",
000081 => x"E8BD8010",
000082 => x"E3A030FF",
000083 => x"E1A03C13",
000084 => x"E1E0E003",
000085 => x"E3E02A0F",
000086 => x"E5123F8F",
000087 => x"E003300E",
000088 => x"E1833C11",
000089 => x"E5023F8F",
000090 => x"E8BD8010",
000091 => x"E20000FF",
000092 => x"E3500007",
000093 => x"E3A02000",
000094 => x"8A00000A",
000095 => x"E2403004",
000096 => x"E3500003",
000097 => x"E20320FF",
000098 => x"9A000005",
000099 => x"E3E03A0F",
000100 => x"E5130F8B",
000101 => x"E1A02182",
000102 => x"E1A00230",
000103 => x"E20000FF",
000104 => x"E1A0F00E",
000105 => x"E1A02180",
000106 => x"E3E03A0F",
000107 => x"E5130F8F",
000108 => x"E1A00230",
000109 => x"E20000FF",
000110 => x"E1A0F00E",
000111 => x"E3E02A0F",
000112 => x"E5123EFB",
000113 => x"E3130002",
000114 => x"E3E00000",
000115 => x"15120EFF",
000116 => x"E1A0F00E",
000117 => x"E3E02A0F",
000118 => x"E5123EFB",
000119 => x"E3130001",
000120 => x"0AFFFFFC",
000121 => x"E20030FF",
000122 => x"E5023EFF",
000123 => x"E1A0F00E",
000124 => x"E20000FF",
000125 => x"E3500001",
000126 => x"E3812B01",
000127 => x"03E03A0F",
000128 => x"E3811B09",
000129 => x"13E03A0F",
000130 => x"05031CFF",
000131 => x"15032CFF",
000132 => x"E1A0F00E",
000133 => x"E3E03A0F",
000134 => x"E5030CFB",
000135 => x"E1A0F00E",
000136 => x"E3E02A0F",
000137 => x"E5123CFF",
000138 => x"E3130C01",
000139 => x"1AFFFFFC",
000140 => x"E5020CEF",
000141 => x"E5123CFF",
000142 => x"E3833C01",
000143 => x"E5023CFF",
000144 => x"E3E02A0F",
000145 => x"E5123CFF",
000146 => x"E3130C01",
000147 => x"1AFFFFFC",
000148 => x"E5120CEF",
000149 => x"E1A0F00E",
000150 => x"E3E01A0F",
000151 => x"E5113CF7",
000152 => x"E20000FF",
000153 => x"E3A02001",
000154 => x"E1833012",
000155 => x"E5013CF7",
000156 => x"E1A0F00E",
000157 => x"E20000FF",
000158 => x"E3A02001",
000159 => x"E1A02012",
000160 => x"E3E01A0F",
000161 => x"E5113CF7",
000162 => x"E1E02002",
000163 => x"E0033002",
000164 => x"E5013CF7",
000165 => x"E1A0F00E",
000166 => x"E3E02A0F",
000167 => x"E5123BE7",
000168 => x"E1A01420",
000169 => x"E3C33080",
000170 => x"E5023BE7",
000171 => x"E5020BEF",
000172 => x"E5021BEB",
000173 => x"E5123BE7",
000174 => x"E3833080",
000175 => x"E5023BE7",
000176 => x"E1A0F00E",
000177 => x"E92D4030",
000178 => x"E3A0C090",
000179 => x"E20140FE",
000180 => x"E3E0EA0F",
000181 => x"E5DD500F",
000182 => x"E20000FF",
000183 => x"E50E4BE3",
000184 => x"E20110FF",
000185 => x"E50ECBFF",
000186 => x"E1A04002",
000187 => x"E203C0FF",
000188 => x"E51E3BFF",
000189 => x"E3130002",
000190 => x"1AFFFFFC",
000191 => x"E51E3BFF",
000192 => x"E3130080",
000193 => x"13E00000",
000194 => x"18BD8030",
000195 => x"E35C0000",
000196 => x"0A000012",
000197 => x"E24C3001",
000198 => x"E203C0FF",
000199 => x"E35C0001",
000200 => x"01A02424",
000201 => x"03E03A0F",
000202 => x"13E03A0F",
000203 => x"05032BE3",
000204 => x"15034BE3",
000205 => x"E3E02A0F",
000206 => x"E3A03010",
000207 => x"E5023BFF",
000208 => x"E5123BFF",
000209 => x"E3130002",
000210 => x"1AFFFFFC",
000211 => x"E5123BFF",
000212 => x"E3130080",
000213 => x"0AFFFFEC",
000214 => x"E3E00001",
000215 => x"E8BD8030",
000216 => x"E3500077",
000217 => x"1A00000C",
000218 => x"E3E03A0F",
000219 => x"E3A02050",
000220 => x"E5035BE3",
000221 => x"E5032BFF",
000222 => x"E1A02003",
000223 => x"E5123BFF",
000224 => x"E3130002",
000225 => x"1AFFFFFC",
000226 => x"E5123BFF",
000227 => x"E2130080",
000228 => x"08BD8030",
000229 => x"E3E00002",
000230 => x"E8BD8030",
000231 => x"E3500072",
000232 => x"13E00003",
000233 => x"18BD8030",
000234 => x"E3813001",
000235 => x"E3E02A0F",
000236 => x"E3A01090",
000237 => x"E5023BE3",
000238 => x"E5021BFF",
000239 => x"E5123BFF",
000240 => x"E3130002",
000241 => x"1AFFFFFC",
000242 => x"E5123BFF",
000243 => x"E3130080",
000244 => x"1AFFFFEF",
000245 => x"E3A03068",
000246 => x"E5023BFF",
000247 => x"E3E00A0F",
000248 => x"E5103BFF",
000249 => x"E3130002",
000250 => x"1AFFFFFC",
000251 => x"E5100BE3",
000252 => x"E8BD8030",
000253 => x"E20000FF",
000254 => x"E350000F",
000255 => x"979FF100",
000256 => x"EA00000F",
000257 => x"000104C4",
000258 => x"000104BC",
000259 => x"000104B4",
000260 => x"000104AC",
000261 => x"000104A4",
000262 => x"0001049C",
000263 => x"00010494",
000264 => x"0001048C",
000265 => x"00010484",
000266 => x"0001047C",
000267 => x"00010474",
000268 => x"0001046C",
000269 => x"00010464",
000270 => x"0001045C",
000271 => x"00010454",
000272 => x"0001044C",
000273 => x"E3A00000",
000274 => x"E1A0F00E",
000275 => x"EE1F0F1F",
000276 => x"E1A0F00E",
000277 => x"EE1E0F1E",
000278 => x"E1A0F00E",
000279 => x"EE1D0F1D",
000280 => x"E1A0F00E",
000281 => x"EE1C0F1C",
000282 => x"E1A0F00E",
000283 => x"EE1B0F1B",
000284 => x"E1A0F00E",
000285 => x"EE1A0F1A",
000286 => x"E1A0F00E",
000287 => x"EE190F19",
000288 => x"E1A0F00E",
000289 => x"EE180F18",
000290 => x"E1A0F00E",
000291 => x"EE170F17",
000292 => x"E1A0F00E",
000293 => x"EE160F16",
000294 => x"E1A0F00E",
000295 => x"EE150F15",
000296 => x"E1A0F00E",
000297 => x"EE140F14",
000298 => x"E1A0F00E",
000299 => x"EE130F13",
000300 => x"E1A0F00E",
000301 => x"EE120F12",
000302 => x"E1A0F00E",
000303 => x"EE110F11",
000304 => x"E1A0F00E",
000305 => x"EE100F10",
000306 => x"E1A0F00E",
000307 => x"E20110FF",
000308 => x"E2411006",
000309 => x"E3510007",
000310 => x"979FF101",
000311 => x"EA000008",
000312 => x"00010508",
000313 => x"00010504",
000314 => x"00010504",
000315 => x"00010504",
000316 => x"00010504",
000317 => x"00010510",
000318 => x"00010518",
000319 => x"00010500",
000320 => x"EE0D0F1D",
000321 => x"E1A0F00E",
000322 => x"EE060F16",
000323 => x"E1A0F00E",
000324 => x"EE0B0F1B",
000325 => x"E1A0F00E",
000326 => x"EE0C0F1C",
000327 => x"E1A0F00E",
000328 => x"E92D4010",
000329 => x"E1A04000",
000330 => x"E5D00000",
000331 => x"E3500000",
000332 => x"1A000003",
000333 => x"EA000005",
000334 => x"E5F40001",
000335 => x"E3500000",
000336 => x"0A000002",
000337 => x"EBFFFF22",
000338 => x"E3500000",
000339 => x"CAFFFFF9",
000340 => x"E1A00004",
000341 => x"E8BD8010",
000342 => x"E92D4070",
000343 => x"E2514000",
000344 => x"E1A05000",
000345 => x"E20260FF",
000346 => x"DA00000B",
000347 => x"EBFFFF12",
000348 => x"E3700001",
000349 => x"E20030FF",
000350 => x"0A000005",
000351 => x"E3560001",
000352 => x"E5C53000",
000353 => x"E1A00003",
000354 => x"E2855001",
000355 => x"0A000005",
000356 => x"E2444001",
000357 => x"E3540000",
000358 => x"CAFFFFF3",
000359 => x"E59F300C",
000360 => x"E5C53000",
000361 => x"E8BD8070",
000362 => x"EBFFFF09",
000363 => x"EAFFFFF7",
000364 => x"000110F4",
000365 => x"E92D4030",
000366 => x"E2514000",
000367 => x"E1A05000",
000368 => x"D8BD8030",
000369 => x"E4D50001",
000370 => x"EBFFFF01",
000371 => x"E2544001",
000372 => x"1AFFFFFB",
000373 => x"E8BD8030",
000374 => x"E92D4010",
000375 => x"E20240FF",
000376 => x"E3540008",
000377 => x"83A04008",
000378 => x"8A000001",
000379 => x"E3540000",
000380 => x"03A04001",
000381 => x"E1A02001",
000382 => x"E1A0E004",
000383 => x"E1A0310E",
000384 => x"E35E0001",
000385 => x"E2433004",
000386 => x"E1A0C000",
000387 => x"81A0C330",
000388 => x"E24E3001",
000389 => x"E20CC00F",
000390 => x"E203E0FF",
000391 => x"E35C0009",
000392 => x"E28C3030",
000393 => x"828C3037",
000394 => x"E35E0000",
000395 => x"E4C23001",
000396 => x"1AFFFFF1",
000397 => x"E2443001",
000398 => x"E20330FF",
000399 => x"E0813003",
000400 => x"E5C3E001",
000401 => x"E8BD8010",
000402 => x"E92D4010",
000403 => x"E1A04000",
000404 => x"E3540007",
000405 => x"E3A01010",
000406 => x"E3A00001",
000407 => x"9A000001",
000408 => x"E3A00000",
000409 => x"E8BD8010",
000410 => x"EBFFFEE0",
000411 => x"E3A00006",
000412 => x"EBFFFEF8",
000413 => x"E3A00000",
000414 => x"EBFFFEE8",
000415 => x"E1A00584",
000416 => x"E8BD4010",
000417 => x"EAFFFEE5",
000418 => x"E0603280",
000419 => x"E0800103",
000420 => x"E0800100",
000421 => x"E1A00200",
000422 => x"E3500000",
000423 => x"D1A0F00E",
000424 => x"E1A00000",
000425 => x"E2500001",
000426 => x"1AFFFFFC",
000427 => x"E1A0F00E",
000428 => x"E212C0FF",
000429 => x"0A00000B",
000430 => x"E5D02000",
000431 => x"E5D13000",
000432 => x"E1520003",
000433 => x"0A000004",
000434 => x"EA000008",
000435 => x"E5F02001",
000436 => x"E5F13001",
000437 => x"E1520003",
000438 => x"1A000004",
000439 => x"E24C3001",
000440 => x"E213C0FF",
000441 => x"1AFFFFF8",
000442 => x"E3A00001",
000443 => x"E1A0F00E",
000444 => x"E3A00000",
000445 => x"E1A0F00E",
000446 => x"E92D4030",
000447 => x"E1A04081",
000448 => x"E3540000",
000449 => x"E1A05000",
000450 => x"D3A00000",
000451 => x"D8BD8030",
000452 => x"E3A00000",
000453 => x"E1A01000",
000454 => x"E7D12005",
000455 => x"E2423030",
000456 => x"E082C200",
000457 => x"E3530009",
000458 => x"E242E041",
000459 => x"924C0030",
000460 => x"9A000007",
000461 => x"E0823200",
000462 => x"E35E0005",
000463 => x"E242C061",
000464 => x"92430037",
000465 => x"9A000002",
000466 => x"E0823200",
000467 => x"E35C0005",
000468 => x"92430057",
000469 => x"E2811001",
000470 => x"E1510004",
000471 => x"1AFFFFED",
000472 => x"E8BD8030",
000473 => x"E5D03003",
000474 => x"E5D02002",
000475 => x"E5D01000",
000476 => x"E1833402",
000477 => x"E5D00001",
000478 => x"E1833C01",
000479 => x"E1830800",
000480 => x"E1A0F00E",
000481 => x"E92D45F0",
000482 => x"E3A00000",
000483 => x"E24DD00C",
000484 => x"EBFFFE53",
000485 => x"E3A0100D",
000486 => x"E3A000C3",
000487 => x"EBFFFF4A",
000488 => x"E3A00063",
000489 => x"EBFFFEBB",
000490 => x"E3A00006",
000491 => x"EBFFFF10",
000492 => x"E3A01006",
000493 => x"E3800008",
000494 => x"EBFFFF43",
000495 => x"E3A0000D",
000496 => x"EBFFFF0B",
000497 => x"E1A008A0",
000498 => x"E1E00000",
000499 => x"E200000F",
000500 => x"E3500001",
000501 => x"03A04030",
000502 => x"028DA007",
000503 => x"0A00001A",
000504 => x"E3500002",
000505 => x"0A000070",
000506 => x"E59F07F8",
000507 => x"EBFFFF4B",
000508 => x"E59F07F4",
000509 => x"EBFFFF49",
000510 => x"E59F07F0",
000511 => x"EBFFFF47",
000512 => x"E59F07EC",
000513 => x"EBFFFF45",
000514 => x"E59F07E8",
000515 => x"EBFFFF43",
000516 => x"E59F07E4",
000517 => x"EBFFFF41",
000518 => x"E59F07E0",
000519 => x"EBFFFF3F",
000520 => x"E59F07DC",
000521 => x"EBFFFF3D",
000522 => x"E59F07D8",
000523 => x"EBFFFF3B",
000524 => x"E59F07D4",
000525 => x"EBFFFF39",
000526 => x"E59F07D0",
000527 => x"EBFFFF37",
000528 => x"E28DA007",
000529 => x"EBFFFE5C",
000530 => x"E1A04000",
000531 => x"E3A0000D",
000532 => x"EBFFFEE7",
000533 => x"E3100801",
000534 => x"03A06001",
000535 => x"03A050A0",
000536 => x"1A000035",
000537 => x"E3A04000",
000538 => x"E59F07A4",
000539 => x"EBFFFF2B",
000540 => x"E1A01005",
000541 => x"E1A02004",
000542 => x"E3A03002",
000543 => x"E3A00072",
000544 => x"E58D4000",
000545 => x"EBFFFE8E",
000546 => x"E1A01005",
000547 => x"E5CD0007",
000548 => x"E3A02001",
000549 => x"E3A03002",
000550 => x"E3A00072",
000551 => x"E58D4000",
000552 => x"EBFFFE87",
000553 => x"E3A02002",
000554 => x"E1A03002",
000555 => x"E5CD0008",
000556 => x"E1A01005",
000557 => x"E3A00072",
000558 => x"E58D4000",
000559 => x"EBFFFE80",
000560 => x"E3A03002",
000561 => x"E5CD0009",
000562 => x"E1A01005",
000563 => x"E3A00072",
000564 => x"E3A02003",
000565 => x"E58D4000",
000566 => x"EBFFFE79",
000567 => x"E5DD3007",
000568 => x"E20000FF",
000569 => x"E3530053",
000570 => x"E5CD000A",
000571 => x"1A000002",
000572 => x"E5DD3008",
000573 => x"E353004D",
000574 => x"0A000062",
000575 => x"E59F0714",
000576 => x"EBFFFF06",
000577 => x"E3560000",
000578 => x"0AFFFFCD",
000579 => x"E59F0708",
000580 => x"EBFFFF02",
000581 => x"E3A0100D",
000582 => x"E3A00000",
000583 => x"EBFFFEEA",
000584 => x"E3A00006",
000585 => x"EBFFFEB2",
000586 => x"E3A01006",
000587 => x"E3C00008",
000588 => x"EBFFFEE5",
000589 => x"E3A0F000",
000590 => x"EAFFFFFE",
000591 => x"E3540034",
000592 => x"0A000028",
000593 => x"CA00001B",
000594 => x"E3540031",
000595 => x"0A000035",
000596 => x"DA000097",
000597 => x"E3540032",
000598 => x"0A0000A1",
000599 => x"E3540033",
000600 => x"1A000097",
000601 => x"E1A00004",
000602 => x"EBFFFE19",
000603 => x"E59F06AC",
000604 => x"EBFFFEEA",
000605 => x"E1A0000A",
000606 => x"E3A01002",
000607 => x"E3A02001",
000608 => x"EBFFFEF4",
000609 => x"E3A01002",
000610 => x"E1A0000A",
000611 => x"EBFFFF59",
000612 => x"E21010FF",
000613 => x"11A05001",
000614 => x"13A06000",
000615 => x"1AFFFFB0",
000616 => x"E59F067C",
000617 => x"EBFFFEDD",
000618 => x"EAFFFFA5",
000619 => x"E3A04033",
000620 => x"E28DA007",
000621 => x"EAFFFFA4",
000622 => x"E3540066",
000623 => x"0A00002A",
000624 => x"DA0000A5",
000625 => x"E3540068",
000626 => x"0A000107",
000627 => x"E3540072",
000628 => x"1A00007B",
000629 => x"E1A00004",
000630 => x"EBFFFDFD",
000631 => x"E3A006FF",
000632 => x"E280F20F",
000633 => x"EAFFFFFE",
000634 => x"E1A00004",
000635 => x"EBFFFDF8",
000636 => x"E59F0628",
000637 => x"EBFFFEC9",
000638 => x"E1A0000A",
000639 => x"E3A01002",
000640 => x"E3A02001",
000641 => x"EBFFFED3",
000642 => x"E1A0000A",
000643 => x"E3A01002",
000644 => x"EBFFFF38",
000645 => x"E21080FF",
000646 => x"1A00009C",
000647 => x"E59F0604",
000648 => x"EBFFFEBE",
000649 => x"EAFFFF86",
000650 => x"E1A00004",
000651 => x"EBFFFDE8",
000652 => x"E59F05F4",
000653 => x"EBFFFEB9",
000654 => x"E1A0000A",
000655 => x"E3A01004",
000656 => x"E3A02000",
000657 => x"EBFFFEC3",
000658 => x"E5DD3007",
000659 => x"E3530053",
000660 => x"1A000002",
000661 => x"E5DD3008",
000662 => x"E353004D",
000663 => x"0A00010D",
000664 => x"E59F05C8",
000665 => x"EBFFFEAD",
000666 => x"EAFFFF75",
000667 => x"E1A00004",
000668 => x"EBFFFDD7",
000669 => x"E59F05B8",
000670 => x"EBFFFEA8",
000671 => x"E59F05B4",
000672 => x"EBFFFEA6",
000673 => x"EAFFFF6E",
000674 => x"E5DD3009",
000675 => x"E3530042",
000676 => x"1AFFFF99",
000677 => x"E3500052",
000678 => x"1AFFFF97",
000679 => x"E1A01005",
000680 => x"E3A02004",
000681 => x"E2433040",
000682 => x"E2800020",
000683 => x"E58D4000",
000684 => x"EBFFFE03",
000685 => x"E1A01005",
000686 => x"E5CD0007",
000687 => x"E3A02005",
000688 => x"E3A03002",
000689 => x"E3A00072",
000690 => x"E58D4000",
000691 => x"EBFFFDFC",
000692 => x"E1A01005",
000693 => x"E5CD0008",
000694 => x"E3A02006",
000695 => x"E3A03002",
000696 => x"E3A00072",
000697 => x"E58D4000",
000698 => x"EBFFFDF5",
000699 => x"E1A01005",
000700 => x"E5CD0009",
000701 => x"E3A02007",
000702 => x"E3A03002",
000703 => x"E3A00072",
000704 => x"E58D4000",
000705 => x"EBFFFDEE",
000706 => x"E5CD000A",
000707 => x"E1A0000A",
000708 => x"EBFFFF13",
000709 => x"E2907004",
000710 => x"0A000022",
000711 => x"E1A06004",
000712 => x"E2842008",
000713 => x"E1A01005",
000714 => x"E3A03002",
000715 => x"E3A00072",
000716 => x"E58D6000",
000717 => x"EBFFFDE2",
000718 => x"E2842009",
000719 => x"E5CD0007",
000720 => x"E1A01005",
000721 => x"E3A03002",
000722 => x"E3A00072",
000723 => x"E58D6000",
000724 => x"EBFFFDDB",
000725 => x"E284200A",
000726 => x"E5CD0008",
000727 => x"E1A01005",
000728 => x"E3A03002",
000729 => x"E3A00072",
000730 => x"E58D6000",
000731 => x"EBFFFDD4",
000732 => x"E284200B",
000733 => x"E5CD0009",
000734 => x"E1A01005",
000735 => x"E3A03002",
000736 => x"E3A00072",
000737 => x"E58D6000",
000738 => x"EBFFFDCD",
000739 => x"E5CD000A",
000740 => x"E1A0000A",
000741 => x"EBFFFEF2",
000742 => x"E4840004",
000743 => x"E1540007",
000744 => x"13540902",
000745 => x"3AFFFFDD",
000746 => x"E59F048C",
000747 => x"EBFFFE5B",
000748 => x"EAFFFF55",
000749 => x"E3740001",
000750 => x"0AFFFF21",
000751 => x"E3540030",
000752 => x"0A000004",
000753 => x"E20400FF",
000754 => x"EBFFFD81",
000755 => x"E59F046C",
000756 => x"EBFFFE52",
000757 => x"EAFFFF1A",
000758 => x"E1A00004",
000759 => x"EBFFFD7C",
000760 => x"EAFFFF49",
000761 => x"E1A00004",
000762 => x"EBFFFD79",
000763 => x"E59F0450",
000764 => x"EBFFFE4A",
000765 => x"EBFFFD70",
000766 => x"E3700001",
000767 => x"0AFFFFFC",
000768 => x"EBFFFD6D",
000769 => x"E3700001",
000770 => x"1AFFFFFC",
000771 => x"E3A05000",
000772 => x"EA000001",
000773 => x"E3550902",
000774 => x"0A00000C",
000775 => x"E5954000",
000776 => x"E1A00C24",
000777 => x"EBFFFD6A",
000778 => x"E1A00824",
000779 => x"EBFFFD68",
000780 => x"E1A00424",
000781 => x"EBFFFD66",
000782 => x"E1A00004",
000783 => x"EBFFFD64",
000784 => x"EBFFFD5D",
000785 => x"E3700001",
000786 => x"E2855004",
000787 => x"0AFFFFF0",
000788 => x"E59F03F0",
000789 => x"EBFFFE31",
000790 => x"EAFFFEF9",
000791 => x"E3540035",
000792 => x"0A0000AC",
000793 => x"E3540061",
000794 => x"1AFFFFD5",
000795 => x"E1A00004",
000796 => x"EBFFFD57",
000797 => x"E59F03D0",
000798 => x"EBFFFE28",
000799 => x"E59F03CC",
000800 => x"EBFFFE26",
000801 => x"E59F03C8",
000802 => x"EBFFFE24",
000803 => x"EAFFFEEC",
000804 => x"E59F03C0",
000805 => x"EBFFFE21",
000806 => x"E1A0000A",
000807 => x"E3A01004",
000808 => x"E3A02000",
000809 => x"EBFFFE2B",
000810 => x"E5DD3007",
000811 => x"E3530053",
000812 => x"1A000002",
000813 => x"E5DD2008",
000814 => x"E352004D",
000815 => x"0A000004",
000816 => x"E59F0394",
000817 => x"EBFFFE15",
000818 => x"E59F0390",
000819 => x"EBFFFE13",
000820 => x"EAFFFEDB",
000821 => x"E5DD1009",
000822 => x"E3510042",
000823 => x"1AFFFFF7",
000824 => x"E5DD000A",
000825 => x"E3500052",
000826 => x"1AFFFFF4",
000827 => x"E3A04000",
000828 => x"E5C43000",
000829 => x"E1A00000",
000830 => x"E5C42001",
000831 => x"E1A00000",
000832 => x"E5C41002",
000833 => x"E1A00000",
000834 => x"E5C40003",
000835 => x"E1A00000",
000836 => x"E241103E",
000837 => x"E1A0000A",
000838 => x"E1A02004",
000839 => x"EBFFFE0D",
000840 => x"E5DD3007",
000841 => x"E5C43004",
000842 => x"E5DD2008",
000843 => x"E5C42005",
000844 => x"E5DD3009",
000845 => x"E5C43006",
000846 => x"E5DD200A",
000847 => x"E1A0000A",
000848 => x"E5C42007",
000849 => x"EBFFFE86",
000850 => x"E3A03CFF",
000851 => x"E28330FC",
000852 => x"E1500003",
000853 => x"E1A05000",
000854 => x"8A000098",
000855 => x"E3700004",
000856 => x"12844008",
000857 => x"1280600B",
000858 => x"0A000006",
000859 => x"EBFFFD12",
000860 => x"E3700001",
000861 => x"0AFFFFFC",
000862 => x"E1560004",
000863 => x"E5C40000",
000864 => x"E2844001",
000865 => x"1AFFFFF8",
000866 => x"E59F02D4",
000867 => x"EBFFFDE3",
000868 => x"E59F02D0",
000869 => x"EBFFFDE1",
000870 => x"E375000C",
000871 => x"0A00000F",
000872 => x"E3A04000",
000873 => x"E285700C",
000874 => x"E1A06004",
000875 => x"E5D45000",
000876 => x"E3A00077",
000877 => x"E1A01008",
000878 => x"E1A02006",
000879 => x"E3A03002",
000880 => x"E58D5000",
000881 => x"EBFFFD3E",
000882 => x"E3500000",
000883 => x"1AFFFFF7",
000884 => x"E2844001",
000885 => x"E1540007",
000886 => x"E1A06004",
000887 => x"1AFFFFF2",
000888 => x"E59F0284",
000889 => x"EBFFFDCD",
000890 => x"EAFFFFB6",
000891 => x"E1A00004",
000892 => x"EBFFFCF7",
000893 => x"E59F0274",
000894 => x"EBFFFDC8",
000895 => x"E59F0270",
000896 => x"EBFFFDC6",
000897 => x"E59F026C",
000898 => x"EBFFFDC4",
000899 => x"E59F0268",
000900 => x"EBFFFDC2",
000901 => x"E59F0264",
000902 => x"EBFFFDC0",
000903 => x"E59F0260",
000904 => x"EBFFFDBE",
000905 => x"E59F025C",
000906 => x"EBFFFDBC",
000907 => x"E59F0258",
000908 => x"EBFFFDBA",
000909 => x"E59F0254",
000910 => x"EBFFFDB8",
000911 => x"E59F0250",
000912 => x"EBFFFDB6",
000913 => x"E59F024C",
000914 => x"EBFFFDB4",
000915 => x"E59F0248",
000916 => x"EBFFFDB2",
000917 => x"E59F0244",
000918 => x"EBFFFDB0",
000919 => x"E59F0240",
000920 => x"EBFFFDAE",
000921 => x"E59F023C",
000922 => x"EBFFFDAC",
000923 => x"E59F0238",
000924 => x"EBFFFDAA",
000925 => x"E59F0234",
000926 => x"EBFFFDA8",
000927 => x"E59F0230",
000928 => x"EBFFFDA6",
000929 => x"E59F022C",
000930 => x"EBFFFDA4",
000931 => x"E59F0228",
000932 => x"EBFFFDA2",
000933 => x"EAFFFE6A",
000934 => x"E5DD3009",
000935 => x"E3530042",
000936 => x"1AFFFEEE",
000937 => x"E5DD300A",
000938 => x"E3530052",
000939 => x"1AFFFEEB",
000940 => x"E3A01004",
000941 => x"E3A02000",
000942 => x"E1A0000A",
000943 => x"EBFFFDA5",
000944 => x"E1A0000A",
000945 => x"EBFFFE26",
000946 => x"E3A03C7F",
000947 => x"E28330F8",
000948 => x"E1500003",
000949 => x"8A000039",
000950 => x"E2905004",
000951 => x"0A000009",
000952 => x"E3A04000",
000953 => x"E3A01004",
000954 => x"E3A02000",
000955 => x"E1A0000A",
000956 => x"EBFFFD98",
000957 => x"E1A0000A",
000958 => x"EBFFFE19",
000959 => x"E4840004",
000960 => x"E1550004",
000961 => x"1AFFFFF6",
000962 => x"E1A00000",
000963 => x"E1A00000",
000964 => x"E1A00000",
000965 => x"EAFFFE7C",
000966 => x"E1A00004",
000967 => x"EBFFFCAC",
000968 => x"E59F0198",
000969 => x"EBFFFD7D",
000970 => x"E1A0000A",
000971 => x"E3A01002",
000972 => x"E3A02001",
000973 => x"EBFFFD87",
000974 => x"E1A0000A",
000975 => x"E3A01002",
000976 => x"EBFFFDEC",
000977 => x"E21060FF",
000978 => x"0AFFFE94",
000979 => x"E59F0170",
000980 => x"EBFFFD72",
000981 => x"E59F016C",
000982 => x"EBFFFD70",
000983 => x"EBFFFC96",
000984 => x"E3700001",
000985 => x"0AFFFFFC",
000986 => x"EBFFFC93",
000987 => x"E3700001",
000988 => x"1AFFFFFC",
000989 => x"E3A05000",
000990 => x"EA000001",
000991 => x"E3540000",
000992 => x"AA000011",
000993 => x"E3A0C000",
000994 => x"E1A02005",
000995 => x"E1A01006",
000996 => x"E3A03002",
000997 => x"E3A00072",
000998 => x"E58DC000",
000999 => x"EBFFFCC8",
001000 => x"E1A04000",
001001 => x"EBFFFC84",
001002 => x"E3700001",
001003 => x"E1A00004",
001004 => x"0AFFFFF1",
001005 => x"E59F0110",
001006 => x"EBFFFD58",
001007 => x"EAFFFF23",
001008 => x"E59F0108",
001009 => x"EBFFFD55",
001010 => x"EAFFFE1D",
001011 => x"EBFFFC80",
001012 => x"E3A03801",
001013 => x"E2855001",
001014 => x"E2433001",
001015 => x"E1550003",
001016 => x"1AFFFFE7",
001017 => x"EAFFFF19",
001018 => x"000110F8",
001019 => x"00011144",
001020 => x"0001118C",
001021 => x"000111D4",
001022 => x"0001121C",
001023 => x"00011264",
001024 => x"000112AC",
001025 => x"00011318",
001026 => x"00011350",
001027 => x"000113B4",
001028 => x"00011418",
001029 => x"000115F0",
001030 => x"00011654",
001031 => x"00011D58",
001032 => x"00011594",
001033 => x"000115D0",
001034 => x"00011680",
001035 => x"00011468",
001036 => x"00011500",
001037 => x"00011CDC",
001038 => x"00011D0C",
001039 => x"00011640",
001040 => x"00011D34",
001041 => x"00011528",
001042 => x"00011570",
001043 => x"00011830",
001044 => x"00011864",
001045 => x"000118D0",
001046 => x"000116A0",
001047 => x"00011748",
001048 => x"00011D28",
001049 => x"00011700",
001050 => x"00011718",
001051 => x"00011738",
001052 => x"00011914",
001053 => x"00011930",
001054 => x"00011950",
001055 => x"00011990",
001056 => x"000119C4",
001057 => x"00011A00",
001058 => x"00011A3C",
001059 => x"00011A60",
001060 => x"00011A9C",
001061 => x"00011AB8",
001062 => x"00011AD0",
001063 => x"00011B18",
001064 => x"00011B58",
001065 => x"00011B90",
001066 => x"00011BB4",
001067 => x"00011BF8",
001068 => x"00011C38",
001069 => x"00011C64",
001070 => x"00011C90",
001071 => x"00011CB4",
001072 => x"0001176C",
001073 => x"000117A8",
001074 => x"000117E8",
001075 => x"00011D7C",
001076 => x"000114DC",
001077 => x"E10F3000",
001078 => x"E3C330C0",
001079 => x"E129F003",
001080 => x"E1A0F00E",
001081 => x"E10F3000",
001082 => x"E38330C0",
001083 => x"E129F003",
001084 => x"E1A0F00E",
001085 => x"00000000",
001086 => x"0D0A0D0A",
001087 => x"0D0A2B2D",
001088 => x"2D2D2D2D",
001089 => x"2D2D2D2D",
001090 => x"2D2D2D2D",
001091 => x"2D2D2D2D",
001092 => x"2D2D2D2D",
001093 => x"2D2D2D2D",
001094 => x"2D2D2D2D",
001095 => x"2D2D2D2D",
001096 => x"2D2D2D2D",
001097 => x"2D2D2D2D",
001098 => x"2D2D2D2D",
001099 => x"2D2D2D2D",
001100 => x"2D2D2D2D",
001101 => x"2D2D2D2D",
001102 => x"2D2D2D2D",
001103 => x"2D2D2D2B",
001104 => x"0D0A0000",
001105 => x"7C202020",
001106 => x"203C3C3C",
001107 => x"2053544F",
001108 => x"524D2043",
001109 => x"6F726520",
001110 => x"50726F63",
001111 => x"6573736F",
001112 => x"72205379",
001113 => x"7374656D",
001114 => x"202D2042",
001115 => x"79205374",
001116 => x"65706861",
001117 => x"6E204E6F",
001118 => x"6C74696E",
001119 => x"67203E3E",
001120 => x"3E202020",
001121 => x"207C0D0A",
001122 => x"00000000",
001123 => x"2B2D2D2D",
001124 => x"2D2D2D2D",
001125 => x"2D2D2D2D",
001126 => x"2D2D2D2D",
001127 => x"2D2D2D2D",
001128 => x"2D2D2D2D",
001129 => x"2D2D2D2D",
001130 => x"2D2D2D2D",
001131 => x"2D2D2D2D",
001132 => x"2D2D2D2D",
001133 => x"2D2D2D2D",
001134 => x"2D2D2D2D",
001135 => x"2D2D2D2D",
001136 => x"2D2D2D2D",
001137 => x"2D2D2D2D",
001138 => x"2D2D2D2D",
001139 => x"2D2B0D0A",
001140 => x"00000000",
001141 => x"7C202020",
001142 => x"20202020",
001143 => x"2020426F",
001144 => x"6F746C6F",
001145 => x"61646572",
001146 => x"20666F72",
001147 => x"2053544F",
001148 => x"524D2053",
001149 => x"6F432020",
001150 => x"20566572",
001151 => x"73696F6E",
001152 => x"3A203230",
001153 => x"31323035",
001154 => x"32342D44",
001155 => x"20202020",
001156 => x"20202020",
001157 => x"207C0D0A",
001158 => x"00000000",
001159 => x"7C202020",
001160 => x"20202020",
001161 => x"20202020",
001162 => x"20202020",
001163 => x"436F6E74",
001164 => x"6163743A",
001165 => x"2073746E",
001166 => x"6F6C7469",
001167 => x"6E674067",
001168 => x"6F6F676C",
001169 => x"656D6169",
001170 => x"6C2E636F",
001171 => x"6D202020",
001172 => x"20202020",
001173 => x"20202020",
001174 => x"20202020",
001175 => x"207C0D0A",
001176 => x"00000000",
001177 => x"2B2D2D2D",
001178 => x"2D2D2D2D",
001179 => x"2D2D2D2D",
001180 => x"2D2D2D2D",
001181 => x"2D2D2D2D",
001182 => x"2D2D2D2D",
001183 => x"2D2D2D2D",
001184 => x"2D2D2D2D",
001185 => x"2D2D2D2D",
001186 => x"2D2D2D2D",
001187 => x"2D2D2D2D",
001188 => x"2D2D2D2D",
001189 => x"2D2D2D2D",
001190 => x"2D2D2D2D",
001191 => x"2D2D2D2D",
001192 => x"2D2D2D2D",
001193 => x"2D2B0D0A",
001194 => x"0D0A0000",
001195 => x"203C2057",
001196 => x"656C636F",
001197 => x"6D652074",
001198 => x"6F207468",
001199 => x"65205354",
001200 => x"4F524D20",
001201 => x"536F4320",
001202 => x"626F6F74",
001203 => x"6C6F6164",
001204 => x"65722063",
001205 => x"6F6E736F",
001206 => x"6C652120",
001207 => x"3E0D0A20",
001208 => x"3C205365",
001209 => x"6C656374",
001210 => x"20616E20",
001211 => x"6F706572",
001212 => x"6174696F",
001213 => x"6E206672",
001214 => x"6F6D2074",
001215 => x"6865206D",
001216 => x"656E7520",
001217 => x"62656C6F",
001218 => x"77206F72",
001219 => x"20707265",
001220 => x"7373203E",
001221 => x"0D0A0000",
001222 => x"203C2074",
001223 => x"68652062",
001224 => x"6F6F7420",
001225 => x"6B657920",
001226 => x"666F7220",
001227 => x"696D6D65",
001228 => x"64696174",
001229 => x"65206170",
001230 => x"706C6963",
001231 => x"6174696F",
001232 => x"6E207374",
001233 => x"6172742E",
001234 => x"203E0D0A",
001235 => x"0D0A0000",
001236 => x"2030202D",
001237 => x"20626F6F",
001238 => x"74206672",
001239 => x"6F6D2063",
001240 => x"6F726520",
001241 => x"52414D20",
001242 => x"28737461",
001243 => x"72742061",
001244 => x"70706C69",
001245 => x"63617469",
001246 => x"6F6E290D",
001247 => x"0A203120",
001248 => x"2D207072",
001249 => x"6F677261",
001250 => x"6D20636F",
001251 => x"72652052",
001252 => x"414D2076",
001253 => x"69612055",
001254 => x"4152545F",
001255 => x"300D0A20",
001256 => x"32202D20",
001257 => x"636F7265",
001258 => x"2052414D",
001259 => x"2064756D",
001260 => x"700D0A00",
001261 => x"2033202D",
001262 => x"20626F6F",
001263 => x"74206672",
001264 => x"6F6D2049",
001265 => x"32432045",
001266 => x"4550524F",
001267 => x"4D0D0A20",
001268 => x"34202D20",
001269 => x"70726F67",
001270 => x"72616D20",
001271 => x"49324320",
001272 => x"45455052",
001273 => x"4F4D2076",
001274 => x"69612055",
001275 => x"4152545F",
001276 => x"300D0A20",
001277 => x"35202D20",
001278 => x"73686F77",
001279 => x"20636F6E",
001280 => x"74656E74",
001281 => x"206F6620",
001282 => x"49324320",
001283 => x"45455052",
001284 => x"4F4D0D0A",
001285 => x"00000000",
001286 => x"2061202D",
001287 => x"20617574",
001288 => x"6F6D6174",
001289 => x"69632062",
001290 => x"6F6F7420",
001291 => x"636F6E66",
001292 => x"69677572",
001293 => x"6174696F",
001294 => x"6E0D0A20",
001295 => x"68202D20",
001296 => x"68656C70",
001297 => x"0D0A2072",
001298 => x"202D2072",
001299 => x"65737461",
001300 => x"72742073",
001301 => x"79737465",
001302 => x"6D0D0A0D",
001303 => x"0A53656C",
001304 => x"6563743A",
001305 => x"20000000",
001306 => x"0D0A0D0A",
001307 => x"4170706C",
001308 => x"69636174",
001309 => x"696F6E20",
001310 => x"77696C6C",
001311 => x"20737461",
001312 => x"72742061",
001313 => x"75746F6D",
001314 => x"61746963",
001315 => x"616C6C79",
001316 => x"20616674",
001317 => x"65722064",
001318 => x"6F776E6C",
001319 => x"6F61642E",
001320 => x"0D0A2D3E",
001321 => x"20576169",
001322 => x"74696E67",
001323 => x"20666F72",
001324 => x"20277374",
001325 => x"6F726D5F",
001326 => x"70726F67",
001327 => x"72616D2E",
001328 => x"62696E27",
001329 => x"20696E20",
001330 => x"62797465",
001331 => x"2D737472",
001332 => x"65616D20",
001333 => x"6D6F6465",
001334 => x"2E2E2E00",
001335 => x"20455252",
001336 => x"4F522120",
001337 => x"50726F67",
001338 => x"72616D20",
001339 => x"66696C65",
001340 => x"20746F6F",
001341 => x"20626967",
001342 => x"210D0A0D",
001343 => x"0A000000",
001344 => x"20496E76",
001345 => x"616C6964",
001346 => x"2070726F",
001347 => x"6772616D",
001348 => x"6D696E67",
001349 => x"2066696C",
001350 => x"65210D0A",
001351 => x"0D0A5365",
001352 => x"6C656374",
001353 => x"3A200000",
001354 => x"0D0A0D0A",
001355 => x"41626F72",
001356 => x"74206475",
001357 => x"6D70696E",
001358 => x"67206279",
001359 => x"20707265",
001360 => x"7373696E",
001361 => x"6720616E",
001362 => x"79206B65",
001363 => x"792E0D0A",
001364 => x"50726573",
001365 => x"7320616E",
001366 => x"79206B65",
001367 => x"7920746F",
001368 => x"20636F6E",
001369 => x"74696E75",
001370 => x"652E0D0A",
001371 => x"0D0A0000",
001372 => x"0D0A0D0A",
001373 => x"44756D70",
001374 => x"696E6720",
001375 => x"636F6D70",
001376 => x"6C657465",
001377 => x"642E0D0A",
001378 => x"0D0A5365",
001379 => x"6C656374",
001380 => x"3A200000",
001381 => x"0D0A0D0A",
001382 => x"456E7465",
001383 => x"72206465",
001384 => x"76696365",
001385 => x"20616464",
001386 => x"72657373",
001387 => x"20283278",
001388 => x"20686578",
001389 => x"5F636861",
001390 => x"72732C20",
001391 => x"73657420",
001392 => x"4C534220",
001393 => x"746F2027",
001394 => x"3027293A",
001395 => x"20000000",
001396 => x"20496E76",
001397 => x"616C6964",
001398 => x"20616464",
001399 => x"72657373",
001400 => x"210D0A0D",
001401 => x"0A53656C",
001402 => x"6563743A",
001403 => x"20000000",
001404 => x"0D0A4170",
001405 => x"706C6963",
001406 => x"6174696F",
001407 => x"6E207769",
001408 => x"6C6C2073",
001409 => x"74617274",
001410 => x"20617574",
001411 => x"6F6D6174",
001412 => x"6963616C",
001413 => x"6C792061",
001414 => x"66746572",
001415 => x"2075706C",
001416 => x"6F61642E",
001417 => x"0D0A2D3E",
001418 => x"204C6F61",
001419 => x"64696E67",
001420 => x"20626F6F",
001421 => x"7420696D",
001422 => x"6167652E",
001423 => x"2E2E0000",
001424 => x"2055706C",
001425 => x"6F616420",
001426 => x"636F6D70",
001427 => x"6C657465",
001428 => x"0D0A0000",
001429 => x"20496E76",
001430 => x"616C6964",
001431 => x"20626F6F",
001432 => x"74206465",
001433 => x"76696365",
001434 => x"206F7220",
001435 => x"66696C65",
001436 => x"210D0A0D",
001437 => x"0A53656C",
001438 => x"6563743A",
001439 => x"20000000",
001440 => x"0D0A496E",
001441 => x"76616C69",
001442 => x"64206164",
001443 => x"64726573",
001444 => x"73210D0A",
001445 => x"0D0A5365",
001446 => x"6C656374",
001447 => x"3A200000",
001448 => x"0D0A4461",
001449 => x"74612077",
001450 => x"696C6C20",
001451 => x"6F766572",
001452 => x"77726974",
001453 => x"65205241",
001454 => x"4D20636F",
001455 => x"6E74656E",
001456 => x"74210D0A",
001457 => x"2D3E2057",
001458 => x"61697469",
001459 => x"6E672066",
001460 => x"6F722027",
001461 => x"73746F72",
001462 => x"6D5F7072",
001463 => x"6F677261",
001464 => x"6D2E6269",
001465 => x"6E272069",
001466 => x"6E206279",
001467 => x"74652D73",
001468 => x"74726561",
001469 => x"6D206D6F",
001470 => x"64652E2E",
001471 => x"2E000000",
001472 => x"20446F77",
001473 => x"6E6C6F61",
001474 => x"6420636F",
001475 => x"6D706C65",
001476 => x"7465640D",
001477 => x"0A000000",
001478 => x"57726974",
001479 => x"696E6720",
001480 => x"62756666",
001481 => x"65722074",
001482 => x"6F206932",
001483 => x"63204545",
001484 => x"50524F4D",
001485 => x"2E2E2E00",
001486 => x"20436F6D",
001487 => x"706C6574",
001488 => x"65640D0A",
001489 => x"0D0A0000",
001490 => x"20496E76",
001491 => x"616C6964",
001492 => x"20626F6F",
001493 => x"74206465",
001494 => x"76696365",
001495 => x"206F7220",
001496 => x"66696C65",
001497 => x"210D0A0D",
001498 => x"0A000000",
001499 => x"0D0A0D0A",
001500 => x"456E7465",
001501 => x"72206465",
001502 => x"76696365",
001503 => x"20616464",
001504 => x"72657373",
001505 => x"20283220",
001506 => x"6865782D",
001507 => x"63686172",
001508 => x"732C2073",
001509 => x"6574204C",
001510 => x"53422074",
001511 => x"6F202730",
001512 => x"27293A20",
001513 => x"00000000",
001514 => x"0D0A0D0A",
001515 => x"41626F72",
001516 => x"74206475",
001517 => x"6D70696E",
001518 => x"67206279",
001519 => x"20707265",
001520 => x"7373696E",
001521 => x"6720616E",
001522 => x"79206B65",
001523 => x"792E2049",
001524 => x"66206E6F",
001525 => x"20646174",
001526 => x"61206973",
001527 => x"2073686F",
001528 => x"776E2C0D",
001529 => x"0A000000",
001530 => x"74686520",
001531 => x"73656C65",
001532 => x"63746564",
001533 => x"20646576",
001534 => x"69636520",
001535 => x"6973206E",
001536 => x"6F742072",
001537 => x"6573706F",
001538 => x"6E64696E",
001539 => x"672E2050",
001540 => x"72657373",
001541 => x"20616E79",
001542 => x"206B6579",
001543 => x"20746F20",
001544 => x"636F6E74",
001545 => x"696E7565",
001546 => x"2E0D0A0D",
001547 => x"0A000000",
001548 => x"0D0A0D0A",
001549 => x"4175746F",
001550 => x"6D617469",
001551 => x"6320626F",
001552 => x"6F742063",
001553 => x"6F6E6669",
001554 => x"67757261",
001555 => x"74696F6E",
001556 => x"20666F72",
001557 => x"20706F77",
001558 => x"65722D75",
001559 => x"703A0D0A",
001560 => x"00000000",
001561 => x"5B333231",
001562 => x"305D2063",
001563 => x"6F6E6669",
001564 => x"67757261",
001565 => x"74696F6E",
001566 => x"20444950",
001567 => x"20737769",
001568 => x"7463680D",
001569 => x"0A203030",
001570 => x"3030202D",
001571 => x"20537461",
001572 => x"72742062",
001573 => x"6F6F746C",
001574 => x"6F616465",
001575 => x"7220636F",
001576 => x"6E736F6C",
001577 => x"650D0A20",
001578 => x"30303031",
001579 => x"202D2041",
001580 => x"75746F6D",
001581 => x"61746963",
001582 => x"20626F6F",
001583 => x"74206672",
001584 => x"6F6D2063",
001585 => x"6F726520",
001586 => x"52414D0D",
001587 => x"0A000000",
001588 => x"20303031",
001589 => x"30202D20",
001590 => x"4175746F",
001591 => x"6D617469",
001592 => x"6320626F",
001593 => x"6F742066",
001594 => x"726F6D20",
001595 => x"49324320",
001596 => x"45455052",
001597 => x"4F4D2028",
001598 => x"41646472",
001599 => x"65737320",
001600 => x"30784130",
001601 => x"290D0A0D",
001602 => x"0A53656C",
001603 => x"6563743A",
001604 => x"20000000",
001605 => x"0D0A0D0A",
001606 => x"53544F52",
001607 => x"4D20536F",
001608 => x"4320626F",
001609 => x"6F746C6F",
001610 => x"61646572",
001611 => x"0D0A0000",
001612 => x"2730273A",
001613 => x"20457865",
001614 => x"63757465",
001615 => x"2070726F",
001616 => x"6772616D",
001617 => x"20696E20",
001618 => x"52414D2E",
001619 => x"0D0A0000",
001620 => x"2731273A",
001621 => x"20577269",
001622 => x"74652027",
001623 => x"73746F72",
001624 => x"6D5F7072",
001625 => x"6F677261",
001626 => x"6D2E6269",
001627 => x"6E272074",
001628 => x"6F207468",
001629 => x"6520636F",
001630 => x"72652773",
001631 => x"2052414D",
001632 => x"20766961",
001633 => x"20554152",
001634 => x"542E0D0A",
001635 => x"00000000",
001636 => x"2732273A",
001637 => x"20507269",
001638 => x"6E742063",
001639 => x"75727265",
001640 => x"6E742063",
001641 => x"6F6E7465",
001642 => x"6E74206F",
001643 => x"6620636F",
001644 => x"6D706C65",
001645 => x"74652063",
001646 => x"6F726520",
001647 => x"52414D2E",
001648 => x"0D0A0000",
001649 => x"2733273A",
001650 => x"204C6F61",
001651 => x"6420626F",
001652 => x"6F742069",
001653 => x"6D616765",
001654 => x"2066726F",
001655 => x"6D204545",
001656 => x"50524F4D",
001657 => x"20616E64",
001658 => x"20737461",
001659 => x"72742061",
001660 => x"70706C69",
001661 => x"63617469",
001662 => x"6F6E2E0D",
001663 => x"0A000000",
001664 => x"2734273A",
001665 => x"20577269",
001666 => x"74652027",
001667 => x"73746F72",
001668 => x"6D5F7072",
001669 => x"6F677261",
001670 => x"6D2E6269",
001671 => x"6E272074",
001672 => x"6F204932",
001673 => x"43204545",
001674 => x"50524F4D",
001675 => x"20766961",
001676 => x"20554152",
001677 => x"542E0D0A",
001678 => x"00000000",
001679 => x"2735273A",
001680 => x"20507269",
001681 => x"6E742063",
001682 => x"6F6E7465",
001683 => x"6E74206F",
001684 => x"66204932",
001685 => x"43204545",
001686 => x"50524F4D",
001687 => x"2E0D0A00",
001688 => x"2761273A",
001689 => x"2053686F",
001690 => x"77204449",
001691 => x"50207377",
001692 => x"69746368",
001693 => x"20636F6E",
001694 => x"66696775",
001695 => x"72617469",
001696 => x"6F6E7320",
001697 => x"666F7220",
001698 => x"6175746F",
001699 => x"6D617469",
001700 => x"6320626F",
001701 => x"6F742E0D",
001702 => x"0A000000",
001703 => x"2768273A",
001704 => x"2053686F",
001705 => x"77207468",
001706 => x"69732073",
001707 => x"63726565",
001708 => x"6E2E0D0A",
001709 => x"00000000",
001710 => x"2772273A",
001711 => x"20526573",
001712 => x"65742073",
001713 => x"79737465",
001714 => x"6D2E0D0A",
001715 => x"0D0A0000",
001716 => x"426F6F74",
001717 => x"20454550",
001718 => x"524F4D3A",
001719 => x"20323478",
001720 => x"786E6E6E",
001721 => x"20286C69",
001722 => x"6B652032",
001723 => x"34414136",
001724 => x"34292C20",
001725 => x"37206269",
001726 => x"74206164",
001727 => x"64726573",
001728 => x"73202B20",
001729 => x"646F6E74",
001730 => x"2D636172",
001731 => x"65206269",
001732 => x"742C0D0A",
001733 => x"00000000",
001734 => x"636F6E6E",
001735 => x"65637465",
001736 => x"6420746F",
001737 => x"20493243",
001738 => x"5F434F4E",
001739 => x"54524F4C",
001740 => x"4C45525F",
001741 => x"302C206F",
001742 => x"70657261",
001743 => x"74696E67",
001744 => x"20667265",
001745 => x"7175656E",
001746 => x"63792069",
001747 => x"73203130",
001748 => x"306B487A",
001749 => x"2C0D0A00",
001750 => x"6D617869",
001751 => x"6D756D20",
001752 => x"45455052",
001753 => x"4F4D2073",
001754 => x"697A6520",
001755 => x"3D203635",
001756 => x"35333620",
001757 => x"62797465",
001758 => x"203D3E20",
001759 => x"31362062",
001760 => x"69742061",
001761 => x"64647265",
001762 => x"73736573",
001763 => x"2C0D0A00",
001764 => x"66697865",
001765 => x"6420626F",
001766 => x"6F742064",
001767 => x"65766963",
001768 => x"65206164",
001769 => x"64726573",
001770 => x"733A2030",
001771 => x"7841300D",
001772 => x"0A0D0A00",
001773 => x"5465726D",
001774 => x"696E616C",
001775 => x"20736574",
001776 => x"75703A20",
001777 => x"39363030",
001778 => x"20626175",
001779 => x"642C2038",
001780 => x"20646174",
001781 => x"61206269",
001782 => x"74732C20",
001783 => x"6E6F2070",
001784 => x"61726974",
001785 => x"792C2031",
001786 => x"2073746F",
001787 => x"70206269",
001788 => x"740D0A0D",
001789 => x"0A000000",
001790 => x"466F7220",
001791 => x"6D6F7265",
001792 => x"20696E66",
001793 => x"6F726D61",
001794 => x"74696F6E",
001795 => x"20736565",
001796 => x"20746865",
001797 => x"2053544F",
001798 => x"524D2043",
001799 => x"6F726520",
001800 => x"2F205354",
001801 => x"4F524D20",
001802 => x"536F4320",
001803 => x"64617461",
001804 => x"73686565",
001805 => x"740D0A00",
001806 => x"68747470",
001807 => x"3A2F2F6F",
001808 => x"70656E63",
001809 => x"6F726573",
001810 => x"2E6F7267",
001811 => x"2F70726F",
001812 => x"6A656374",
001813 => x"2C73746F",
001814 => x"726D5F63",
001815 => x"6F72650D",
001816 => x"0A000000",
001817 => x"68747470",
001818 => x"3A2F2F6F",
001819 => x"70656E63",
001820 => x"6F726573",
001821 => x"2E6F7267",
001822 => x"2F70726F",
001823 => x"6A656374",
001824 => x"2C73746F",
001825 => x"726D5F73",
001826 => x"6F630D0A",
001827 => x"00000000",
001828 => x"436F6E74",
001829 => x"6163743A",
001830 => x"2073746E",
001831 => x"6F6C7469",
001832 => x"6E674067",
001833 => x"6F6F676C",
001834 => x"656D6169",
001835 => x"6C2E636F",
001836 => x"6D0D0A00",
001837 => x"28632920",
001838 => x"32303132",
001839 => x"20627920",
001840 => x"53746570",
001841 => x"68616E20",
001842 => x"4E6F6C74",
001843 => x"696E670D",
001844 => x"0A0D0A53",
001845 => x"656C6563",
001846 => x"743A2000",
001847 => x"0D0A0D0A",
001848 => x"5765276C",
001849 => x"6C207365",
001850 => x"6E642079",
001851 => x"6F752062",
001852 => x"61636B20",
001853 => x"2D20746F",
001854 => x"20746865",
001855 => x"20667574",
001856 => x"75726521",
001857 => x"2E0D0A0D",
001858 => x"0A000000",
001859 => x"202D2044",
001860 => x"6F63746F",
001861 => x"7220456D",
001862 => x"6D657420",
001863 => x"4C2E2042",
001864 => x"726F776E",
001865 => x"0D0A0D0A",
001866 => x"53656C65",
001867 => x"63743A20",
001868 => x"00000000",
001869 => x"20496E76",
001870 => x"616C6964",
001871 => x"206F7065",
001872 => x"72617469",
001873 => x"6F6E210D",
001874 => x"0A547279",
001875 => x"20616761",
001876 => x"696E3A20",
001877 => x"00000000",
001878 => x"0D0A0D0A",
001879 => x"2D3E2053",
001880 => x"74617274",
001881 => x"696E6720",
001882 => x"6170706C",
001883 => x"69636174",
001884 => x"696F6E2E",
001885 => x"2E2E0D0A",
001886 => x"0D0A0000",
001887 => x"0D0A0D0A",
001888 => x"41626F72",
001889 => x"74656421",
001890 => x"00000000",
others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;